`default_nettype none

module static_arbiter_16 (input wire clock, message_interface_nonblocking.producer out0, message_interface_nonblocking.producer out1, message_interface_nonblocking.producer out2, message_interface_nonblocking.producer out3, message_interface_nonblocking.producer out4, message_interface_nonblocking.producer out5, message_interface_nonblocking.producer out6, message_interface_nonblocking.producer out7, message_interface_nonblocking.producer out8, message_interface_nonblocking.producer out9, message_interface_nonblocking.producer out10, message_interface_nonblocking.producer out11, message_interface_nonblocking.producer out12, message_interface_nonblocking.producer out13, message_interface_nonblocking.producer out14, message_interface_nonblocking.producer out15, message_interface.consumer in0, message_interface.consumer in1, message_interface.consumer in2, message_interface.consumer in3, message_interface.consumer in4, message_interface.consumer in5, message_interface.consumer in6, message_interface.consumer in7, message_interface.consumer in8, message_interface.consumer in9, message_interface.consumer in10, message_interface.consumer in11, message_interface.consumer in12, message_interface.consumer in13, message_interface.consumer in14, message_interface.consumer in15);
  wire [16-1:0] req [16-1:0];
  wire [16-1:0] req_prefix [16-1:0];
  wire [16-1:0] ack [16-1:0];
  wire [16-1:0] any_ack;
  
parPrefix2OR_16 req_prefix_tree_0 (.in(req[0]),.out(req_prefix[0]));
parPrefix2OR_16 req_prefix_tree_1 (.in(req[1]),.out(req_prefix[1]));
parPrefix2OR_16 req_prefix_tree_2 (.in(req[2]),.out(req_prefix[2]));
parPrefix2OR_16 req_prefix_tree_3 (.in(req[3]),.out(req_prefix[3]));
parPrefix2OR_16 req_prefix_tree_4 (.in(req[4]),.out(req_prefix[4]));
parPrefix2OR_16 req_prefix_tree_5 (.in(req[5]),.out(req_prefix[5]));
parPrefix2OR_16 req_prefix_tree_6 (.in(req[6]),.out(req_prefix[6]));
parPrefix2OR_16 req_prefix_tree_7 (.in(req[7]),.out(req_prefix[7]));
parPrefix2OR_16 req_prefix_tree_8 (.in(req[8]),.out(req_prefix[8]));
parPrefix2OR_16 req_prefix_tree_9 (.in(req[9]),.out(req_prefix[9]));
parPrefix2OR_16 req_prefix_tree_10 (.in(req[10]),.out(req_prefix[10]));
parPrefix2OR_16 req_prefix_tree_11 (.in(req[11]),.out(req_prefix[11]));
parPrefix2OR_16 req_prefix_tree_12 (.in(req[12]),.out(req_prefix[12]));
parPrefix2OR_16 req_prefix_tree_13 (.in(req[13]),.out(req_prefix[13]));
parPrefix2OR_16 req_prefix_tree_14 (.in(req[14]),.out(req_prefix[14]));
parPrefix2OR_16 req_prefix_tree_15 (.in(req[15]),.out(req_prefix[15]));
  assign req[0][0] = in0.valid && (in0.to == 0);
  assign ack[0][0] = req[0][0];
  assign req[1][0] = in0.valid && (in0.to == 1);
  assign ack[0][1] = req[1][0];
  assign req[2][0] = in0.valid && (in0.to == 2);
  assign ack[0][2] = req[2][0];
  assign req[3][0] = in0.valid && (in0.to == 3);
  assign ack[0][3] = req[3][0];
  assign req[4][0] = in0.valid && (in0.to == 4);
  assign ack[0][4] = req[4][0];
  assign req[5][0] = in0.valid && (in0.to == 5);
  assign ack[0][5] = req[5][0];
  assign req[6][0] = in0.valid && (in0.to == 6);
  assign ack[0][6] = req[6][0];
  assign req[7][0] = in0.valid && (in0.to == 7);
  assign ack[0][7] = req[7][0];
  assign req[8][0] = in0.valid && (in0.to == 8);
  assign ack[0][8] = req[8][0];
  assign req[9][0] = in0.valid && (in0.to == 9);
  assign ack[0][9] = req[9][0];
  assign req[10][0] = in0.valid && (in0.to == 10);
  assign ack[0][10] = req[10][0];
  assign req[11][0] = in0.valid && (in0.to == 11);
  assign ack[0][11] = req[11][0];
  assign req[12][0] = in0.valid && (in0.to == 12);
  assign ack[0][12] = req[12][0];
  assign req[13][0] = in0.valid && (in0.to == 13);
  assign ack[0][13] = req[13][0];
  assign req[14][0] = in0.valid && (in0.to == 14);
  assign ack[0][14] = req[14][0];
  assign req[15][0] = in0.valid && (in0.to == 15);
  assign ack[0][15] = req[15][0];
  assign any_ack[0] = ack[0][0]||ack[0][1]||ack[0][2]||ack[0][3]||ack[0][4]||ack[0][5]||ack[0][6]||ack[0][7]||ack[0][8]||ack[0][9]||ack[0][10]||ack[0][11]||ack[0][12]||ack[0][13]||ack[0][14]||ack[0][15];
  assign in0.ack = any_ack[0];
  assign out0.valid = any_ack[0];
  assign out0.to = any_ack[0] ? in0.to : 0;
  assign out0.from = any_ack[0] ? in0.from : 0;
  assign out0.data = any_ack[0] ? in0.data : 0;
  assign req[0][1] = in1.valid && (in1.to == 0);
  assign ack[1][0] = req[0][1] && !req_prefix[0][1-1];
  assign req[1][1] = in1.valid && (in1.to == 1);
  assign ack[1][1] = req[1][1] && !req_prefix[1][1-1];
  assign req[2][1] = in1.valid && (in1.to == 2);
  assign ack[1][2] = req[2][1] && !req_prefix[2][1-1];
  assign req[3][1] = in1.valid && (in1.to == 3);
  assign ack[1][3] = req[3][1] && !req_prefix[3][1-1];
  assign req[4][1] = in1.valid && (in1.to == 4);
  assign ack[1][4] = req[4][1] && !req_prefix[4][1-1];
  assign req[5][1] = in1.valid && (in1.to == 5);
  assign ack[1][5] = req[5][1] && !req_prefix[5][1-1];
  assign req[6][1] = in1.valid && (in1.to == 6);
  assign ack[1][6] = req[6][1] && !req_prefix[6][1-1];
  assign req[7][1] = in1.valid && (in1.to == 7);
  assign ack[1][7] = req[7][1] && !req_prefix[7][1-1];
  assign req[8][1] = in1.valid && (in1.to == 8);
  assign ack[1][8] = req[8][1] && !req_prefix[8][1-1];
  assign req[9][1] = in1.valid && (in1.to == 9);
  assign ack[1][9] = req[9][1] && !req_prefix[9][1-1];
  assign req[10][1] = in1.valid && (in1.to == 10);
  assign ack[1][10] = req[10][1] && !req_prefix[10][1-1];
  assign req[11][1] = in1.valid && (in1.to == 11);
  assign ack[1][11] = req[11][1] && !req_prefix[11][1-1];
  assign req[12][1] = in1.valid && (in1.to == 12);
  assign ack[1][12] = req[12][1] && !req_prefix[12][1-1];
  assign req[13][1] = in1.valid && (in1.to == 13);
  assign ack[1][13] = req[13][1] && !req_prefix[13][1-1];
  assign req[14][1] = in1.valid && (in1.to == 14);
  assign ack[1][14] = req[14][1] && !req_prefix[14][1-1];
  assign req[15][1] = in1.valid && (in1.to == 15);
  assign ack[1][15] = req[15][1] && !req_prefix[15][1-1];
  assign any_ack[1] = ack[1][0]||ack[1][1]||ack[1][2]||ack[1][3]||ack[1][4]||ack[1][5]||ack[1][6]||ack[1][7]||ack[1][8]||ack[1][9]||ack[1][10]||ack[1][11]||ack[1][12]||ack[1][13]||ack[1][14]||ack[1][15];
  assign in1.ack = any_ack[1];
  assign out1.valid = any_ack[1];
  assign out1.to = any_ack[1] ? in1.to : 0;
  assign out1.from = any_ack[1] ? in1.from : 0;
  assign out1.data = any_ack[1] ? in1.data : 0;
  assign req[0][2] = in2.valid && (in2.to == 0);
  assign ack[2][0] = req[0][2] && !req_prefix[0][2-1];
  assign req[1][2] = in2.valid && (in2.to == 1);
  assign ack[2][1] = req[1][2] && !req_prefix[1][2-1];
  assign req[2][2] = in2.valid && (in2.to == 2);
  assign ack[2][2] = req[2][2] && !req_prefix[2][2-1];
  assign req[3][2] = in2.valid && (in2.to == 3);
  assign ack[2][3] = req[3][2] && !req_prefix[3][2-1];
  assign req[4][2] = in2.valid && (in2.to == 4);
  assign ack[2][4] = req[4][2] && !req_prefix[4][2-1];
  assign req[5][2] = in2.valid && (in2.to == 5);
  assign ack[2][5] = req[5][2] && !req_prefix[5][2-1];
  assign req[6][2] = in2.valid && (in2.to == 6);
  assign ack[2][6] = req[6][2] && !req_prefix[6][2-1];
  assign req[7][2] = in2.valid && (in2.to == 7);
  assign ack[2][7] = req[7][2] && !req_prefix[7][2-1];
  assign req[8][2] = in2.valid && (in2.to == 8);
  assign ack[2][8] = req[8][2] && !req_prefix[8][2-1];
  assign req[9][2] = in2.valid && (in2.to == 9);
  assign ack[2][9] = req[9][2] && !req_prefix[9][2-1];
  assign req[10][2] = in2.valid && (in2.to == 10);
  assign ack[2][10] = req[10][2] && !req_prefix[10][2-1];
  assign req[11][2] = in2.valid && (in2.to == 11);
  assign ack[2][11] = req[11][2] && !req_prefix[11][2-1];
  assign req[12][2] = in2.valid && (in2.to == 12);
  assign ack[2][12] = req[12][2] && !req_prefix[12][2-1];
  assign req[13][2] = in2.valid && (in2.to == 13);
  assign ack[2][13] = req[13][2] && !req_prefix[13][2-1];
  assign req[14][2] = in2.valid && (in2.to == 14);
  assign ack[2][14] = req[14][2] && !req_prefix[14][2-1];
  assign req[15][2] = in2.valid && (in2.to == 15);
  assign ack[2][15] = req[15][2] && !req_prefix[15][2-1];
  assign any_ack[2] = ack[2][0]||ack[2][1]||ack[2][2]||ack[2][3]||ack[2][4]||ack[2][5]||ack[2][6]||ack[2][7]||ack[2][8]||ack[2][9]||ack[2][10]||ack[2][11]||ack[2][12]||ack[2][13]||ack[2][14]||ack[2][15];
  assign in2.ack = any_ack[2];
  assign out2.valid = any_ack[2];
  assign out2.to = any_ack[2] ? in2.to : 0;
  assign out2.from = any_ack[2] ? in2.from : 0;
  assign out2.data = any_ack[2] ? in2.data : 0;
  assign req[0][3] = in3.valid && (in3.to == 0);
  assign ack[3][0] = req[0][3] && !req_prefix[0][3-1];
  assign req[1][3] = in3.valid && (in3.to == 1);
  assign ack[3][1] = req[1][3] && !req_prefix[1][3-1];
  assign req[2][3] = in3.valid && (in3.to == 2);
  assign ack[3][2] = req[2][3] && !req_prefix[2][3-1];
  assign req[3][3] = in3.valid && (in3.to == 3);
  assign ack[3][3] = req[3][3] && !req_prefix[3][3-1];
  assign req[4][3] = in3.valid && (in3.to == 4);
  assign ack[3][4] = req[4][3] && !req_prefix[4][3-1];
  assign req[5][3] = in3.valid && (in3.to == 5);
  assign ack[3][5] = req[5][3] && !req_prefix[5][3-1];
  assign req[6][3] = in3.valid && (in3.to == 6);
  assign ack[3][6] = req[6][3] && !req_prefix[6][3-1];
  assign req[7][3] = in3.valid && (in3.to == 7);
  assign ack[3][7] = req[7][3] && !req_prefix[7][3-1];
  assign req[8][3] = in3.valid && (in3.to == 8);
  assign ack[3][8] = req[8][3] && !req_prefix[8][3-1];
  assign req[9][3] = in3.valid && (in3.to == 9);
  assign ack[3][9] = req[9][3] && !req_prefix[9][3-1];
  assign req[10][3] = in3.valid && (in3.to == 10);
  assign ack[3][10] = req[10][3] && !req_prefix[10][3-1];
  assign req[11][3] = in3.valid && (in3.to == 11);
  assign ack[3][11] = req[11][3] && !req_prefix[11][3-1];
  assign req[12][3] = in3.valid && (in3.to == 12);
  assign ack[3][12] = req[12][3] && !req_prefix[12][3-1];
  assign req[13][3] = in3.valid && (in3.to == 13);
  assign ack[3][13] = req[13][3] && !req_prefix[13][3-1];
  assign req[14][3] = in3.valid && (in3.to == 14);
  assign ack[3][14] = req[14][3] && !req_prefix[14][3-1];
  assign req[15][3] = in3.valid && (in3.to == 15);
  assign ack[3][15] = req[15][3] && !req_prefix[15][3-1];
  assign any_ack[3] = ack[3][0]||ack[3][1]||ack[3][2]||ack[3][3]||ack[3][4]||ack[3][5]||ack[3][6]||ack[3][7]||ack[3][8]||ack[3][9]||ack[3][10]||ack[3][11]||ack[3][12]||ack[3][13]||ack[3][14]||ack[3][15];
  assign in3.ack = any_ack[3];
  assign out3.valid = any_ack[3];
  assign out3.to = any_ack[3] ? in3.to : 0;
  assign out3.from = any_ack[3] ? in3.from : 0;
  assign out3.data = any_ack[3] ? in3.data : 0;
  assign req[0][4] = in4.valid && (in4.to == 0);
  assign ack[4][0] = req[0][4] && !req_prefix[0][4-1];
  assign req[1][4] = in4.valid && (in4.to == 1);
  assign ack[4][1] = req[1][4] && !req_prefix[1][4-1];
  assign req[2][4] = in4.valid && (in4.to == 2);
  assign ack[4][2] = req[2][4] && !req_prefix[2][4-1];
  assign req[3][4] = in4.valid && (in4.to == 3);
  assign ack[4][3] = req[3][4] && !req_prefix[3][4-1];
  assign req[4][4] = in4.valid && (in4.to == 4);
  assign ack[4][4] = req[4][4] && !req_prefix[4][4-1];
  assign req[5][4] = in4.valid && (in4.to == 5);
  assign ack[4][5] = req[5][4] && !req_prefix[5][4-1];
  assign req[6][4] = in4.valid && (in4.to == 6);
  assign ack[4][6] = req[6][4] && !req_prefix[6][4-1];
  assign req[7][4] = in4.valid && (in4.to == 7);
  assign ack[4][7] = req[7][4] && !req_prefix[7][4-1];
  assign req[8][4] = in4.valid && (in4.to == 8);
  assign ack[4][8] = req[8][4] && !req_prefix[8][4-1];
  assign req[9][4] = in4.valid && (in4.to == 9);
  assign ack[4][9] = req[9][4] && !req_prefix[9][4-1];
  assign req[10][4] = in4.valid && (in4.to == 10);
  assign ack[4][10] = req[10][4] && !req_prefix[10][4-1];
  assign req[11][4] = in4.valid && (in4.to == 11);
  assign ack[4][11] = req[11][4] && !req_prefix[11][4-1];
  assign req[12][4] = in4.valid && (in4.to == 12);
  assign ack[4][12] = req[12][4] && !req_prefix[12][4-1];
  assign req[13][4] = in4.valid && (in4.to == 13);
  assign ack[4][13] = req[13][4] && !req_prefix[13][4-1];
  assign req[14][4] = in4.valid && (in4.to == 14);
  assign ack[4][14] = req[14][4] && !req_prefix[14][4-1];
  assign req[15][4] = in4.valid && (in4.to == 15);
  assign ack[4][15] = req[15][4] && !req_prefix[15][4-1];
  assign any_ack[4] = ack[4][0]||ack[4][1]||ack[4][2]||ack[4][3]||ack[4][4]||ack[4][5]||ack[4][6]||ack[4][7]||ack[4][8]||ack[4][9]||ack[4][10]||ack[4][11]||ack[4][12]||ack[4][13]||ack[4][14]||ack[4][15];
  assign in4.ack = any_ack[4];
  assign out4.valid = any_ack[4];
  assign out4.to = any_ack[4] ? in4.to : 0;
  assign out4.from = any_ack[4] ? in4.from : 0;
  assign out4.data = any_ack[4] ? in4.data : 0;
  assign req[0][5] = in5.valid && (in5.to == 0);
  assign ack[5][0] = req[0][5] && !req_prefix[0][5-1];
  assign req[1][5] = in5.valid && (in5.to == 1);
  assign ack[5][1] = req[1][5] && !req_prefix[1][5-1];
  assign req[2][5] = in5.valid && (in5.to == 2);
  assign ack[5][2] = req[2][5] && !req_prefix[2][5-1];
  assign req[3][5] = in5.valid && (in5.to == 3);
  assign ack[5][3] = req[3][5] && !req_prefix[3][5-1];
  assign req[4][5] = in5.valid && (in5.to == 4);
  assign ack[5][4] = req[4][5] && !req_prefix[4][5-1];
  assign req[5][5] = in5.valid && (in5.to == 5);
  assign ack[5][5] = req[5][5] && !req_prefix[5][5-1];
  assign req[6][5] = in5.valid && (in5.to == 6);
  assign ack[5][6] = req[6][5] && !req_prefix[6][5-1];
  assign req[7][5] = in5.valid && (in5.to == 7);
  assign ack[5][7] = req[7][5] && !req_prefix[7][5-1];
  assign req[8][5] = in5.valid && (in5.to == 8);
  assign ack[5][8] = req[8][5] && !req_prefix[8][5-1];
  assign req[9][5] = in5.valid && (in5.to == 9);
  assign ack[5][9] = req[9][5] && !req_prefix[9][5-1];
  assign req[10][5] = in5.valid && (in5.to == 10);
  assign ack[5][10] = req[10][5] && !req_prefix[10][5-1];
  assign req[11][5] = in5.valid && (in5.to == 11);
  assign ack[5][11] = req[11][5] && !req_prefix[11][5-1];
  assign req[12][5] = in5.valid && (in5.to == 12);
  assign ack[5][12] = req[12][5] && !req_prefix[12][5-1];
  assign req[13][5] = in5.valid && (in5.to == 13);
  assign ack[5][13] = req[13][5] && !req_prefix[13][5-1];
  assign req[14][5] = in5.valid && (in5.to == 14);
  assign ack[5][14] = req[14][5] && !req_prefix[14][5-1];
  assign req[15][5] = in5.valid && (in5.to == 15);
  assign ack[5][15] = req[15][5] && !req_prefix[15][5-1];
  assign any_ack[5] = ack[5][0]||ack[5][1]||ack[5][2]||ack[5][3]||ack[5][4]||ack[5][5]||ack[5][6]||ack[5][7]||ack[5][8]||ack[5][9]||ack[5][10]||ack[5][11]||ack[5][12]||ack[5][13]||ack[5][14]||ack[5][15];
  assign in5.ack = any_ack[5];
  assign out5.valid = any_ack[5];
  assign out5.to = any_ack[5] ? in5.to : 0;
  assign out5.from = any_ack[5] ? in5.from : 0;
  assign out5.data = any_ack[5] ? in5.data : 0;
  assign req[0][6] = in6.valid && (in6.to == 0);
  assign ack[6][0] = req[0][6] && !req_prefix[0][6-1];
  assign req[1][6] = in6.valid && (in6.to == 1);
  assign ack[6][1] = req[1][6] && !req_prefix[1][6-1];
  assign req[2][6] = in6.valid && (in6.to == 2);
  assign ack[6][2] = req[2][6] && !req_prefix[2][6-1];
  assign req[3][6] = in6.valid && (in6.to == 3);
  assign ack[6][3] = req[3][6] && !req_prefix[3][6-1];
  assign req[4][6] = in6.valid && (in6.to == 4);
  assign ack[6][4] = req[4][6] && !req_prefix[4][6-1];
  assign req[5][6] = in6.valid && (in6.to == 5);
  assign ack[6][5] = req[5][6] && !req_prefix[5][6-1];
  assign req[6][6] = in6.valid && (in6.to == 6);
  assign ack[6][6] = req[6][6] && !req_prefix[6][6-1];
  assign req[7][6] = in6.valid && (in6.to == 7);
  assign ack[6][7] = req[7][6] && !req_prefix[7][6-1];
  assign req[8][6] = in6.valid && (in6.to == 8);
  assign ack[6][8] = req[8][6] && !req_prefix[8][6-1];
  assign req[9][6] = in6.valid && (in6.to == 9);
  assign ack[6][9] = req[9][6] && !req_prefix[9][6-1];
  assign req[10][6] = in6.valid && (in6.to == 10);
  assign ack[6][10] = req[10][6] && !req_prefix[10][6-1];
  assign req[11][6] = in6.valid && (in6.to == 11);
  assign ack[6][11] = req[11][6] && !req_prefix[11][6-1];
  assign req[12][6] = in6.valid && (in6.to == 12);
  assign ack[6][12] = req[12][6] && !req_prefix[12][6-1];
  assign req[13][6] = in6.valid && (in6.to == 13);
  assign ack[6][13] = req[13][6] && !req_prefix[13][6-1];
  assign req[14][6] = in6.valid && (in6.to == 14);
  assign ack[6][14] = req[14][6] && !req_prefix[14][6-1];
  assign req[15][6] = in6.valid && (in6.to == 15);
  assign ack[6][15] = req[15][6] && !req_prefix[15][6-1];
  assign any_ack[6] = ack[6][0]||ack[6][1]||ack[6][2]||ack[6][3]||ack[6][4]||ack[6][5]||ack[6][6]||ack[6][7]||ack[6][8]||ack[6][9]||ack[6][10]||ack[6][11]||ack[6][12]||ack[6][13]||ack[6][14]||ack[6][15];
  assign in6.ack = any_ack[6];
  assign out6.valid = any_ack[6];
  assign out6.to = any_ack[6] ? in6.to : 0;
  assign out6.from = any_ack[6] ? in6.from : 0;
  assign out6.data = any_ack[6] ? in6.data : 0;
  assign req[0][7] = in7.valid && (in7.to == 0);
  assign ack[7][0] = req[0][7] && !req_prefix[0][7-1];
  assign req[1][7] = in7.valid && (in7.to == 1);
  assign ack[7][1] = req[1][7] && !req_prefix[1][7-1];
  assign req[2][7] = in7.valid && (in7.to == 2);
  assign ack[7][2] = req[2][7] && !req_prefix[2][7-1];
  assign req[3][7] = in7.valid && (in7.to == 3);
  assign ack[7][3] = req[3][7] && !req_prefix[3][7-1];
  assign req[4][7] = in7.valid && (in7.to == 4);
  assign ack[7][4] = req[4][7] && !req_prefix[4][7-1];
  assign req[5][7] = in7.valid && (in7.to == 5);
  assign ack[7][5] = req[5][7] && !req_prefix[5][7-1];
  assign req[6][7] = in7.valid && (in7.to == 6);
  assign ack[7][6] = req[6][7] && !req_prefix[6][7-1];
  assign req[7][7] = in7.valid && (in7.to == 7);
  assign ack[7][7] = req[7][7] && !req_prefix[7][7-1];
  assign req[8][7] = in7.valid && (in7.to == 8);
  assign ack[7][8] = req[8][7] && !req_prefix[8][7-1];
  assign req[9][7] = in7.valid && (in7.to == 9);
  assign ack[7][9] = req[9][7] && !req_prefix[9][7-1];
  assign req[10][7] = in7.valid && (in7.to == 10);
  assign ack[7][10] = req[10][7] && !req_prefix[10][7-1];
  assign req[11][7] = in7.valid && (in7.to == 11);
  assign ack[7][11] = req[11][7] && !req_prefix[11][7-1];
  assign req[12][7] = in7.valid && (in7.to == 12);
  assign ack[7][12] = req[12][7] && !req_prefix[12][7-1];
  assign req[13][7] = in7.valid && (in7.to == 13);
  assign ack[7][13] = req[13][7] && !req_prefix[13][7-1];
  assign req[14][7] = in7.valid && (in7.to == 14);
  assign ack[7][14] = req[14][7] && !req_prefix[14][7-1];
  assign req[15][7] = in7.valid && (in7.to == 15);
  assign ack[7][15] = req[15][7] && !req_prefix[15][7-1];
  assign any_ack[7] = ack[7][0]||ack[7][1]||ack[7][2]||ack[7][3]||ack[7][4]||ack[7][5]||ack[7][6]||ack[7][7]||ack[7][8]||ack[7][9]||ack[7][10]||ack[7][11]||ack[7][12]||ack[7][13]||ack[7][14]||ack[7][15];
  assign in7.ack = any_ack[7];
  assign out7.valid = any_ack[7];
  assign out7.to = any_ack[7] ? in7.to : 0;
  assign out7.from = any_ack[7] ? in7.from : 0;
  assign out7.data = any_ack[7] ? in7.data : 0;
  assign req[0][8] = in8.valid && (in8.to == 0);
  assign ack[8][0] = req[0][8] && !req_prefix[0][8-1];
  assign req[1][8] = in8.valid && (in8.to == 1);
  assign ack[8][1] = req[1][8] && !req_prefix[1][8-1];
  assign req[2][8] = in8.valid && (in8.to == 2);
  assign ack[8][2] = req[2][8] && !req_prefix[2][8-1];
  assign req[3][8] = in8.valid && (in8.to == 3);
  assign ack[8][3] = req[3][8] && !req_prefix[3][8-1];
  assign req[4][8] = in8.valid && (in8.to == 4);
  assign ack[8][4] = req[4][8] && !req_prefix[4][8-1];
  assign req[5][8] = in8.valid && (in8.to == 5);
  assign ack[8][5] = req[5][8] && !req_prefix[5][8-1];
  assign req[6][8] = in8.valid && (in8.to == 6);
  assign ack[8][6] = req[6][8] && !req_prefix[6][8-1];
  assign req[7][8] = in8.valid && (in8.to == 7);
  assign ack[8][7] = req[7][8] && !req_prefix[7][8-1];
  assign req[8][8] = in8.valid && (in8.to == 8);
  assign ack[8][8] = req[8][8] && !req_prefix[8][8-1];
  assign req[9][8] = in8.valid && (in8.to == 9);
  assign ack[8][9] = req[9][8] && !req_prefix[9][8-1];
  assign req[10][8] = in8.valid && (in8.to == 10);
  assign ack[8][10] = req[10][8] && !req_prefix[10][8-1];
  assign req[11][8] = in8.valid && (in8.to == 11);
  assign ack[8][11] = req[11][8] && !req_prefix[11][8-1];
  assign req[12][8] = in8.valid && (in8.to == 12);
  assign ack[8][12] = req[12][8] && !req_prefix[12][8-1];
  assign req[13][8] = in8.valid && (in8.to == 13);
  assign ack[8][13] = req[13][8] && !req_prefix[13][8-1];
  assign req[14][8] = in8.valid && (in8.to == 14);
  assign ack[8][14] = req[14][8] && !req_prefix[14][8-1];
  assign req[15][8] = in8.valid && (in8.to == 15);
  assign ack[8][15] = req[15][8] && !req_prefix[15][8-1];
  assign any_ack[8] = ack[8][0]||ack[8][1]||ack[8][2]||ack[8][3]||ack[8][4]||ack[8][5]||ack[8][6]||ack[8][7]||ack[8][8]||ack[8][9]||ack[8][10]||ack[8][11]||ack[8][12]||ack[8][13]||ack[8][14]||ack[8][15];
  assign in8.ack = any_ack[8];
  assign out8.valid = any_ack[8];
  assign out8.to = any_ack[8] ? in8.to : 0;
  assign out8.from = any_ack[8] ? in8.from : 0;
  assign out8.data = any_ack[8] ? in8.data : 0;
  assign req[0][9] = in9.valid && (in9.to == 0);
  assign ack[9][0] = req[0][9] && !req_prefix[0][9-1];
  assign req[1][9] = in9.valid && (in9.to == 1);
  assign ack[9][1] = req[1][9] && !req_prefix[1][9-1];
  assign req[2][9] = in9.valid && (in9.to == 2);
  assign ack[9][2] = req[2][9] && !req_prefix[2][9-1];
  assign req[3][9] = in9.valid && (in9.to == 3);
  assign ack[9][3] = req[3][9] && !req_prefix[3][9-1];
  assign req[4][9] = in9.valid && (in9.to == 4);
  assign ack[9][4] = req[4][9] && !req_prefix[4][9-1];
  assign req[5][9] = in9.valid && (in9.to == 5);
  assign ack[9][5] = req[5][9] && !req_prefix[5][9-1];
  assign req[6][9] = in9.valid && (in9.to == 6);
  assign ack[9][6] = req[6][9] && !req_prefix[6][9-1];
  assign req[7][9] = in9.valid && (in9.to == 7);
  assign ack[9][7] = req[7][9] && !req_prefix[7][9-1];
  assign req[8][9] = in9.valid && (in9.to == 8);
  assign ack[9][8] = req[8][9] && !req_prefix[8][9-1];
  assign req[9][9] = in9.valid && (in9.to == 9);
  assign ack[9][9] = req[9][9] && !req_prefix[9][9-1];
  assign req[10][9] = in9.valid && (in9.to == 10);
  assign ack[9][10] = req[10][9] && !req_prefix[10][9-1];
  assign req[11][9] = in9.valid && (in9.to == 11);
  assign ack[9][11] = req[11][9] && !req_prefix[11][9-1];
  assign req[12][9] = in9.valid && (in9.to == 12);
  assign ack[9][12] = req[12][9] && !req_prefix[12][9-1];
  assign req[13][9] = in9.valid && (in9.to == 13);
  assign ack[9][13] = req[13][9] && !req_prefix[13][9-1];
  assign req[14][9] = in9.valid && (in9.to == 14);
  assign ack[9][14] = req[14][9] && !req_prefix[14][9-1];
  assign req[15][9] = in9.valid && (in9.to == 15);
  assign ack[9][15] = req[15][9] && !req_prefix[15][9-1];
  assign any_ack[9] = ack[9][0]||ack[9][1]||ack[9][2]||ack[9][3]||ack[9][4]||ack[9][5]||ack[9][6]||ack[9][7]||ack[9][8]||ack[9][9]||ack[9][10]||ack[9][11]||ack[9][12]||ack[9][13]||ack[9][14]||ack[9][15];
  assign in9.ack = any_ack[9];
  assign out9.valid = any_ack[9];
  assign out9.to = any_ack[9] ? in9.to : 0;
  assign out9.from = any_ack[9] ? in9.from : 0;
  assign out9.data = any_ack[9] ? in9.data : 0;
  assign req[0][10] = in10.valid && (in10.to == 0);
  assign ack[10][0] = req[0][10] && !req_prefix[0][10-1];
  assign req[1][10] = in10.valid && (in10.to == 1);
  assign ack[10][1] = req[1][10] && !req_prefix[1][10-1];
  assign req[2][10] = in10.valid && (in10.to == 2);
  assign ack[10][2] = req[2][10] && !req_prefix[2][10-1];
  assign req[3][10] = in10.valid && (in10.to == 3);
  assign ack[10][3] = req[3][10] && !req_prefix[3][10-1];
  assign req[4][10] = in10.valid && (in10.to == 4);
  assign ack[10][4] = req[4][10] && !req_prefix[4][10-1];
  assign req[5][10] = in10.valid && (in10.to == 5);
  assign ack[10][5] = req[5][10] && !req_prefix[5][10-1];
  assign req[6][10] = in10.valid && (in10.to == 6);
  assign ack[10][6] = req[6][10] && !req_prefix[6][10-1];
  assign req[7][10] = in10.valid && (in10.to == 7);
  assign ack[10][7] = req[7][10] && !req_prefix[7][10-1];
  assign req[8][10] = in10.valid && (in10.to == 8);
  assign ack[10][8] = req[8][10] && !req_prefix[8][10-1];
  assign req[9][10] = in10.valid && (in10.to == 9);
  assign ack[10][9] = req[9][10] && !req_prefix[9][10-1];
  assign req[10][10] = in10.valid && (in10.to == 10);
  assign ack[10][10] = req[10][10] && !req_prefix[10][10-1];
  assign req[11][10] = in10.valid && (in10.to == 11);
  assign ack[10][11] = req[11][10] && !req_prefix[11][10-1];
  assign req[12][10] = in10.valid && (in10.to == 12);
  assign ack[10][12] = req[12][10] && !req_prefix[12][10-1];
  assign req[13][10] = in10.valid && (in10.to == 13);
  assign ack[10][13] = req[13][10] && !req_prefix[13][10-1];
  assign req[14][10] = in10.valid && (in10.to == 14);
  assign ack[10][14] = req[14][10] && !req_prefix[14][10-1];
  assign req[15][10] = in10.valid && (in10.to == 15);
  assign ack[10][15] = req[15][10] && !req_prefix[15][10-1];
  assign any_ack[10] = ack[10][0]||ack[10][1]||ack[10][2]||ack[10][3]||ack[10][4]||ack[10][5]||ack[10][6]||ack[10][7]||ack[10][8]||ack[10][9]||ack[10][10]||ack[10][11]||ack[10][12]||ack[10][13]||ack[10][14]||ack[10][15];
  assign in10.ack = any_ack[10];
  assign out10.valid = any_ack[10];
  assign out10.to = any_ack[10] ? in10.to : 0;
  assign out10.from = any_ack[10] ? in10.from : 0;
  assign out10.data = any_ack[10] ? in10.data : 0;
  assign req[0][11] = in11.valid && (in11.to == 0);
  assign ack[11][0] = req[0][11] && !req_prefix[0][11-1];
  assign req[1][11] = in11.valid && (in11.to == 1);
  assign ack[11][1] = req[1][11] && !req_prefix[1][11-1];
  assign req[2][11] = in11.valid && (in11.to == 2);
  assign ack[11][2] = req[2][11] && !req_prefix[2][11-1];
  assign req[3][11] = in11.valid && (in11.to == 3);
  assign ack[11][3] = req[3][11] && !req_prefix[3][11-1];
  assign req[4][11] = in11.valid && (in11.to == 4);
  assign ack[11][4] = req[4][11] && !req_prefix[4][11-1];
  assign req[5][11] = in11.valid && (in11.to == 5);
  assign ack[11][5] = req[5][11] && !req_prefix[5][11-1];
  assign req[6][11] = in11.valid && (in11.to == 6);
  assign ack[11][6] = req[6][11] && !req_prefix[6][11-1];
  assign req[7][11] = in11.valid && (in11.to == 7);
  assign ack[11][7] = req[7][11] && !req_prefix[7][11-1];
  assign req[8][11] = in11.valid && (in11.to == 8);
  assign ack[11][8] = req[8][11] && !req_prefix[8][11-1];
  assign req[9][11] = in11.valid && (in11.to == 9);
  assign ack[11][9] = req[9][11] && !req_prefix[9][11-1];
  assign req[10][11] = in11.valid && (in11.to == 10);
  assign ack[11][10] = req[10][11] && !req_prefix[10][11-1];
  assign req[11][11] = in11.valid && (in11.to == 11);
  assign ack[11][11] = req[11][11] && !req_prefix[11][11-1];
  assign req[12][11] = in11.valid && (in11.to == 12);
  assign ack[11][12] = req[12][11] && !req_prefix[12][11-1];
  assign req[13][11] = in11.valid && (in11.to == 13);
  assign ack[11][13] = req[13][11] && !req_prefix[13][11-1];
  assign req[14][11] = in11.valid && (in11.to == 14);
  assign ack[11][14] = req[14][11] && !req_prefix[14][11-1];
  assign req[15][11] = in11.valid && (in11.to == 15);
  assign ack[11][15] = req[15][11] && !req_prefix[15][11-1];
  assign any_ack[11] = ack[11][0]||ack[11][1]||ack[11][2]||ack[11][3]||ack[11][4]||ack[11][5]||ack[11][6]||ack[11][7]||ack[11][8]||ack[11][9]||ack[11][10]||ack[11][11]||ack[11][12]||ack[11][13]||ack[11][14]||ack[11][15];
  assign in11.ack = any_ack[11];
  assign out11.valid = any_ack[11];
  assign out11.to = any_ack[11] ? in11.to : 0;
  assign out11.from = any_ack[11] ? in11.from : 0;
  assign out11.data = any_ack[11] ? in11.data : 0;
  assign req[0][12] = in12.valid && (in12.to == 0);
  assign ack[12][0] = req[0][12] && !req_prefix[0][12-1];
  assign req[1][12] = in12.valid && (in12.to == 1);
  assign ack[12][1] = req[1][12] && !req_prefix[1][12-1];
  assign req[2][12] = in12.valid && (in12.to == 2);
  assign ack[12][2] = req[2][12] && !req_prefix[2][12-1];
  assign req[3][12] = in12.valid && (in12.to == 3);
  assign ack[12][3] = req[3][12] && !req_prefix[3][12-1];
  assign req[4][12] = in12.valid && (in12.to == 4);
  assign ack[12][4] = req[4][12] && !req_prefix[4][12-1];
  assign req[5][12] = in12.valid && (in12.to == 5);
  assign ack[12][5] = req[5][12] && !req_prefix[5][12-1];
  assign req[6][12] = in12.valid && (in12.to == 6);
  assign ack[12][6] = req[6][12] && !req_prefix[6][12-1];
  assign req[7][12] = in12.valid && (in12.to == 7);
  assign ack[12][7] = req[7][12] && !req_prefix[7][12-1];
  assign req[8][12] = in12.valid && (in12.to == 8);
  assign ack[12][8] = req[8][12] && !req_prefix[8][12-1];
  assign req[9][12] = in12.valid && (in12.to == 9);
  assign ack[12][9] = req[9][12] && !req_prefix[9][12-1];
  assign req[10][12] = in12.valid && (in12.to == 10);
  assign ack[12][10] = req[10][12] && !req_prefix[10][12-1];
  assign req[11][12] = in12.valid && (in12.to == 11);
  assign ack[12][11] = req[11][12] && !req_prefix[11][12-1];
  assign req[12][12] = in12.valid && (in12.to == 12);
  assign ack[12][12] = req[12][12] && !req_prefix[12][12-1];
  assign req[13][12] = in12.valid && (in12.to == 13);
  assign ack[12][13] = req[13][12] && !req_prefix[13][12-1];
  assign req[14][12] = in12.valid && (in12.to == 14);
  assign ack[12][14] = req[14][12] && !req_prefix[14][12-1];
  assign req[15][12] = in12.valid && (in12.to == 15);
  assign ack[12][15] = req[15][12] && !req_prefix[15][12-1];
  assign any_ack[12] = ack[12][0]||ack[12][1]||ack[12][2]||ack[12][3]||ack[12][4]||ack[12][5]||ack[12][6]||ack[12][7]||ack[12][8]||ack[12][9]||ack[12][10]||ack[12][11]||ack[12][12]||ack[12][13]||ack[12][14]||ack[12][15];
  assign in12.ack = any_ack[12];
  assign out12.valid = any_ack[12];
  assign out12.to = any_ack[12] ? in12.to : 0;
  assign out12.from = any_ack[12] ? in12.from : 0;
  assign out12.data = any_ack[12] ? in12.data : 0;
  assign req[0][13] = in13.valid && (in13.to == 0);
  assign ack[13][0] = req[0][13] && !req_prefix[0][13-1];
  assign req[1][13] = in13.valid && (in13.to == 1);
  assign ack[13][1] = req[1][13] && !req_prefix[1][13-1];
  assign req[2][13] = in13.valid && (in13.to == 2);
  assign ack[13][2] = req[2][13] && !req_prefix[2][13-1];
  assign req[3][13] = in13.valid && (in13.to == 3);
  assign ack[13][3] = req[3][13] && !req_prefix[3][13-1];
  assign req[4][13] = in13.valid && (in13.to == 4);
  assign ack[13][4] = req[4][13] && !req_prefix[4][13-1];
  assign req[5][13] = in13.valid && (in13.to == 5);
  assign ack[13][5] = req[5][13] && !req_prefix[5][13-1];
  assign req[6][13] = in13.valid && (in13.to == 6);
  assign ack[13][6] = req[6][13] && !req_prefix[6][13-1];
  assign req[7][13] = in13.valid && (in13.to == 7);
  assign ack[13][7] = req[7][13] && !req_prefix[7][13-1];
  assign req[8][13] = in13.valid && (in13.to == 8);
  assign ack[13][8] = req[8][13] && !req_prefix[8][13-1];
  assign req[9][13] = in13.valid && (in13.to == 9);
  assign ack[13][9] = req[9][13] && !req_prefix[9][13-1];
  assign req[10][13] = in13.valid && (in13.to == 10);
  assign ack[13][10] = req[10][13] && !req_prefix[10][13-1];
  assign req[11][13] = in13.valid && (in13.to == 11);
  assign ack[13][11] = req[11][13] && !req_prefix[11][13-1];
  assign req[12][13] = in13.valid && (in13.to == 12);
  assign ack[13][12] = req[12][13] && !req_prefix[12][13-1];
  assign req[13][13] = in13.valid && (in13.to == 13);
  assign ack[13][13] = req[13][13] && !req_prefix[13][13-1];
  assign req[14][13] = in13.valid && (in13.to == 14);
  assign ack[13][14] = req[14][13] && !req_prefix[14][13-1];
  assign req[15][13] = in13.valid && (in13.to == 15);
  assign ack[13][15] = req[15][13] && !req_prefix[15][13-1];
  assign any_ack[13] = ack[13][0]||ack[13][1]||ack[13][2]||ack[13][3]||ack[13][4]||ack[13][5]||ack[13][6]||ack[13][7]||ack[13][8]||ack[13][9]||ack[13][10]||ack[13][11]||ack[13][12]||ack[13][13]||ack[13][14]||ack[13][15];
  assign in13.ack = any_ack[13];
  assign out13.valid = any_ack[13];
  assign out13.to = any_ack[13] ? in13.to : 0;
  assign out13.from = any_ack[13] ? in13.from : 0;
  assign out13.data = any_ack[13] ? in13.data : 0;
  assign req[0][14] = in14.valid && (in14.to == 0);
  assign ack[14][0] = req[0][14] && !req_prefix[0][14-1];
  assign req[1][14] = in14.valid && (in14.to == 1);
  assign ack[14][1] = req[1][14] && !req_prefix[1][14-1];
  assign req[2][14] = in14.valid && (in14.to == 2);
  assign ack[14][2] = req[2][14] && !req_prefix[2][14-1];
  assign req[3][14] = in14.valid && (in14.to == 3);
  assign ack[14][3] = req[3][14] && !req_prefix[3][14-1];
  assign req[4][14] = in14.valid && (in14.to == 4);
  assign ack[14][4] = req[4][14] && !req_prefix[4][14-1];
  assign req[5][14] = in14.valid && (in14.to == 5);
  assign ack[14][5] = req[5][14] && !req_prefix[5][14-1];
  assign req[6][14] = in14.valid && (in14.to == 6);
  assign ack[14][6] = req[6][14] && !req_prefix[6][14-1];
  assign req[7][14] = in14.valid && (in14.to == 7);
  assign ack[14][7] = req[7][14] && !req_prefix[7][14-1];
  assign req[8][14] = in14.valid && (in14.to == 8);
  assign ack[14][8] = req[8][14] && !req_prefix[8][14-1];
  assign req[9][14] = in14.valid && (in14.to == 9);
  assign ack[14][9] = req[9][14] && !req_prefix[9][14-1];
  assign req[10][14] = in14.valid && (in14.to == 10);
  assign ack[14][10] = req[10][14] && !req_prefix[10][14-1];
  assign req[11][14] = in14.valid && (in14.to == 11);
  assign ack[14][11] = req[11][14] && !req_prefix[11][14-1];
  assign req[12][14] = in14.valid && (in14.to == 12);
  assign ack[14][12] = req[12][14] && !req_prefix[12][14-1];
  assign req[13][14] = in14.valid && (in14.to == 13);
  assign ack[14][13] = req[13][14] && !req_prefix[13][14-1];
  assign req[14][14] = in14.valid && (in14.to == 14);
  assign ack[14][14] = req[14][14] && !req_prefix[14][14-1];
  assign req[15][14] = in14.valid && (in14.to == 15);
  assign ack[14][15] = req[15][14] && !req_prefix[15][14-1];
  assign any_ack[14] = ack[14][0]||ack[14][1]||ack[14][2]||ack[14][3]||ack[14][4]||ack[14][5]||ack[14][6]||ack[14][7]||ack[14][8]||ack[14][9]||ack[14][10]||ack[14][11]||ack[14][12]||ack[14][13]||ack[14][14]||ack[14][15];
  assign in14.ack = any_ack[14];
  assign out14.valid = any_ack[14];
  assign out14.to = any_ack[14] ? in14.to : 0;
  assign out14.from = any_ack[14] ? in14.from : 0;
  assign out14.data = any_ack[14] ? in14.data : 0;
  assign req[0][15] = in15.valid && (in15.to == 0);
  assign ack[15][0] = req[0][15] && !req_prefix[0][15-1];
  assign req[1][15] = in15.valid && (in15.to == 1);
  assign ack[15][1] = req[1][15] && !req_prefix[1][15-1];
  assign req[2][15] = in15.valid && (in15.to == 2);
  assign ack[15][2] = req[2][15] && !req_prefix[2][15-1];
  assign req[3][15] = in15.valid && (in15.to == 3);
  assign ack[15][3] = req[3][15] && !req_prefix[3][15-1];
  assign req[4][15] = in15.valid && (in15.to == 4);
  assign ack[15][4] = req[4][15] && !req_prefix[4][15-1];
  assign req[5][15] = in15.valid && (in15.to == 5);
  assign ack[15][5] = req[5][15] && !req_prefix[5][15-1];
  assign req[6][15] = in15.valid && (in15.to == 6);
  assign ack[15][6] = req[6][15] && !req_prefix[6][15-1];
  assign req[7][15] = in15.valid && (in15.to == 7);
  assign ack[15][7] = req[7][15] && !req_prefix[7][15-1];
  assign req[8][15] = in15.valid && (in15.to == 8);
  assign ack[15][8] = req[8][15] && !req_prefix[8][15-1];
  assign req[9][15] = in15.valid && (in15.to == 9);
  assign ack[15][9] = req[9][15] && !req_prefix[9][15-1];
  assign req[10][15] = in15.valid && (in15.to == 10);
  assign ack[15][10] = req[10][15] && !req_prefix[10][15-1];
  assign req[11][15] = in15.valid && (in15.to == 11);
  assign ack[15][11] = req[11][15] && !req_prefix[11][15-1];
  assign req[12][15] = in15.valid && (in15.to == 12);
  assign ack[15][12] = req[12][15] && !req_prefix[12][15-1];
  assign req[13][15] = in15.valid && (in15.to == 13);
  assign ack[15][13] = req[13][15] && !req_prefix[13][15-1];
  assign req[14][15] = in15.valid && (in15.to == 14);
  assign ack[15][14] = req[14][15] && !req_prefix[14][15-1];
  assign req[15][15] = in15.valid && (in15.to == 15);
  assign ack[15][15] = req[15][15] && !req_prefix[15][15-1];
  assign any_ack[15] = ack[15][0]||ack[15][1]||ack[15][2]||ack[15][3]||ack[15][4]||ack[15][5]||ack[15][6]||ack[15][7]||ack[15][8]||ack[15][9]||ack[15][10]||ack[15][11]||ack[15][12]||ack[15][13]||ack[15][14]||ack[15][15];
  assign in15.ack = any_ack[15];
  assign out15.valid = any_ack[15];
  assign out15.to = any_ack[15] ? in15.to : 0;
  assign out15.from = any_ack[15] ? in15.from : 0;
  assign out15.data = any_ack[15] ? in15.data : 0;
`ifdef FORMAL
  // Preconditions:
  correct_from: assume property ((!in0.valid || (in0.from == 0)) && (!in1.valid || (in1.from == 1)) && (!in2.valid || (in2.from == 2)) && (!in3.valid || (in3.from == 3)) && (!in4.valid || (in4.from == 4)) && (!in5.valid || (in5.from == 5)) && (!in6.valid || (in6.from == 6)) && (!in7.valid || (in7.from == 7)) && (!in8.valid || (in8.from == 8)) && (!in9.valid || (in9.from == 9)) && (!in10.valid || (in10.from == 10)) && (!in11.valid || (in11.from == 11)) && (!in12.valid || (in12.from == 12)) && (!in13.valid || (in13.from == 13)) && (!in14.valid || (in14.from == 14)) && (!in15.valid || (in15.from == 15)));
  correct_dest: assume property ((!in0.valid || (in0.to < 16)) && (!in1.valid || (in1.to < 16)) && (!in2.valid || (in2.to < 16)) && (!in3.valid || (in3.to < 16)) && (!in4.valid || (in4.to < 16)) && (!in5.valid || (in5.to < 16)) && (!in6.valid || (in6.to < 16)) && (!in7.valid || (in7.to < 16)) && (!in8.valid || (in8.to < 16)) && (!in9.valid || (in9.to < 16)) && (!in10.valid || (in10.to < 16)) && (!in11.valid || (in11.to < 16)) && (!in12.valid || (in12.to < 16)) && (!in13.valid || (in13.to < 16)) && (!in14.valid || (in14.to < 16)) && (!in15.valid || (in15.to < 16)));
  // Sanity check:
  all_outputs_valid: cover  property (out0.valid && out1.valid && out2.valid && out3.valid && out4.valid && out5.valid && out6.valid && out7.valid && out8.valid && out9.valid && out10.valid && out11.valid && out12.valid && out13.valid && out14.valid && out15.valid);
  // Goals of implementation:
  unique_destination_output: assert property ((!(out0.valid && out1.valid) || (out0.to != out1.to)) && (!(out0.valid && out2.valid) || (out0.to != out2.to)) && (!(out0.valid && out3.valid) || (out0.to != out3.to)) && (!(out0.valid && out4.valid) || (out0.to != out4.to)) && (!(out0.valid && out5.valid) || (out0.to != out5.to)) && (!(out0.valid && out6.valid) || (out0.to != out6.to)) && (!(out0.valid && out7.valid) || (out0.to != out7.to)) && (!(out0.valid && out8.valid) || (out0.to != out8.to)) && (!(out0.valid && out9.valid) || (out0.to != out9.to)) && (!(out0.valid && out10.valid) || (out0.to != out10.to)) && (!(out0.valid && out11.valid) || (out0.to != out11.to)) && (!(out0.valid && out12.valid) || (out0.to != out12.to)) && (!(out0.valid && out13.valid) || (out0.to != out13.to)) && (!(out0.valid && out14.valid) || (out0.to != out14.to)) && (!(out0.valid && out15.valid) || (out0.to != out15.to)) && (!(out1.valid && out0.valid) || (out1.to != out0.to)) && (!(out1.valid && out2.valid) || (out1.to != out2.to)) && (!(out1.valid && out3.valid) || (out1.to != out3.to)) && (!(out1.valid && out4.valid) || (out1.to != out4.to)) && (!(out1.valid && out5.valid) || (out1.to != out5.to)) && (!(out1.valid && out6.valid) || (out1.to != out6.to)) && (!(out1.valid && out7.valid) || (out1.to != out7.to)) && (!(out1.valid && out8.valid) || (out1.to != out8.to)) && (!(out1.valid && out9.valid) || (out1.to != out9.to)) && (!(out1.valid && out10.valid) || (out1.to != out10.to)) && (!(out1.valid && out11.valid) || (out1.to != out11.to)) && (!(out1.valid && out12.valid) || (out1.to != out12.to)) && (!(out1.valid && out13.valid) || (out1.to != out13.to)) && (!(out1.valid && out14.valid) || (out1.to != out14.to)) && (!(out1.valid && out15.valid) || (out1.to != out15.to)) && (!(out2.valid && out0.valid) || (out2.to != out0.to)) && (!(out2.valid && out1.valid) || (out2.to != out1.to)) && (!(out2.valid && out3.valid) || (out2.to != out3.to)) && (!(out2.valid && out4.valid) || (out2.to != out4.to)) && (!(out2.valid && out5.valid) || (out2.to != out5.to)) && (!(out2.valid && out6.valid) || (out2.to != out6.to)) && (!(out2.valid && out7.valid) || (out2.to != out7.to)) && (!(out2.valid && out8.valid) || (out2.to != out8.to)) && (!(out2.valid && out9.valid) || (out2.to != out9.to)) && (!(out2.valid && out10.valid) || (out2.to != out10.to)) && (!(out2.valid && out11.valid) || (out2.to != out11.to)) && (!(out2.valid && out12.valid) || (out2.to != out12.to)) && (!(out2.valid && out13.valid) || (out2.to != out13.to)) && (!(out2.valid && out14.valid) || (out2.to != out14.to)) && (!(out2.valid && out15.valid) || (out2.to != out15.to)) && (!(out3.valid && out0.valid) || (out3.to != out0.to)) && (!(out3.valid && out1.valid) || (out3.to != out1.to)) && (!(out3.valid && out2.valid) || (out3.to != out2.to)) && (!(out3.valid && out4.valid) || (out3.to != out4.to)) && (!(out3.valid && out5.valid) || (out3.to != out5.to)) && (!(out3.valid && out6.valid) || (out3.to != out6.to)) && (!(out3.valid && out7.valid) || (out3.to != out7.to)) && (!(out3.valid && out8.valid) || (out3.to != out8.to)) && (!(out3.valid && out9.valid) || (out3.to != out9.to)) && (!(out3.valid && out10.valid) || (out3.to != out10.to)) && (!(out3.valid && out11.valid) || (out3.to != out11.to)) && (!(out3.valid && out12.valid) || (out3.to != out12.to)) && (!(out3.valid && out13.valid) || (out3.to != out13.to)) && (!(out3.valid && out14.valid) || (out3.to != out14.to)) && (!(out3.valid && out15.valid) || (out3.to != out15.to)) && (!(out4.valid && out0.valid) || (out4.to != out0.to)) && (!(out4.valid && out1.valid) || (out4.to != out1.to)) && (!(out4.valid && out2.valid) || (out4.to != out2.to)) && (!(out4.valid && out3.valid) || (out4.to != out3.to)) && (!(out4.valid && out5.valid) || (out4.to != out5.to)) && (!(out4.valid && out6.valid) || (out4.to != out6.to)) && (!(out4.valid && out7.valid) || (out4.to != out7.to)) && (!(out4.valid && out8.valid) || (out4.to != out8.to)) && (!(out4.valid && out9.valid) || (out4.to != out9.to)) && (!(out4.valid && out10.valid) || (out4.to != out10.to)) && (!(out4.valid && out11.valid) || (out4.to != out11.to)) && (!(out4.valid && out12.valid) || (out4.to != out12.to)) && (!(out4.valid && out13.valid) || (out4.to != out13.to)) && (!(out4.valid && out14.valid) || (out4.to != out14.to)) && (!(out4.valid && out15.valid) || (out4.to != out15.to)) && (!(out5.valid && out0.valid) || (out5.to != out0.to)) && (!(out5.valid && out1.valid) || (out5.to != out1.to)) && (!(out5.valid && out2.valid) || (out5.to != out2.to)) && (!(out5.valid && out3.valid) || (out5.to != out3.to)) && (!(out5.valid && out4.valid) || (out5.to != out4.to)) && (!(out5.valid && out6.valid) || (out5.to != out6.to)) && (!(out5.valid && out7.valid) || (out5.to != out7.to)) && (!(out5.valid && out8.valid) || (out5.to != out8.to)) && (!(out5.valid && out9.valid) || (out5.to != out9.to)) && (!(out5.valid && out10.valid) || (out5.to != out10.to)) && (!(out5.valid && out11.valid) || (out5.to != out11.to)) && (!(out5.valid && out12.valid) || (out5.to != out12.to)) && (!(out5.valid && out13.valid) || (out5.to != out13.to)) && (!(out5.valid && out14.valid) || (out5.to != out14.to)) && (!(out5.valid && out15.valid) || (out5.to != out15.to)) && (!(out6.valid && out0.valid) || (out6.to != out0.to)) && (!(out6.valid && out1.valid) || (out6.to != out1.to)) && (!(out6.valid && out2.valid) || (out6.to != out2.to)) && (!(out6.valid && out3.valid) || (out6.to != out3.to)) && (!(out6.valid && out4.valid) || (out6.to != out4.to)) && (!(out6.valid && out5.valid) || (out6.to != out5.to)) && (!(out6.valid && out7.valid) || (out6.to != out7.to)) && (!(out6.valid && out8.valid) || (out6.to != out8.to)) && (!(out6.valid && out9.valid) || (out6.to != out9.to)) && (!(out6.valid && out10.valid) || (out6.to != out10.to)) && (!(out6.valid && out11.valid) || (out6.to != out11.to)) && (!(out6.valid && out12.valid) || (out6.to != out12.to)) && (!(out6.valid && out13.valid) || (out6.to != out13.to)) && (!(out6.valid && out14.valid) || (out6.to != out14.to)) && (!(out6.valid && out15.valid) || (out6.to != out15.to)) && (!(out7.valid && out0.valid) || (out7.to != out0.to)) && (!(out7.valid && out1.valid) || (out7.to != out1.to)) && (!(out7.valid && out2.valid) || (out7.to != out2.to)) && (!(out7.valid && out3.valid) || (out7.to != out3.to)) && (!(out7.valid && out4.valid) || (out7.to != out4.to)) && (!(out7.valid && out5.valid) || (out7.to != out5.to)) && (!(out7.valid && out6.valid) || (out7.to != out6.to)) && (!(out7.valid && out8.valid) || (out7.to != out8.to)) && (!(out7.valid && out9.valid) || (out7.to != out9.to)) && (!(out7.valid && out10.valid) || (out7.to != out10.to)) && (!(out7.valid && out11.valid) || (out7.to != out11.to)) && (!(out7.valid && out12.valid) || (out7.to != out12.to)) && (!(out7.valid && out13.valid) || (out7.to != out13.to)) && (!(out7.valid && out14.valid) || (out7.to != out14.to)) && (!(out7.valid && out15.valid) || (out7.to != out15.to)) && (!(out8.valid && out0.valid) || (out8.to != out0.to)) && (!(out8.valid && out1.valid) || (out8.to != out1.to)) && (!(out8.valid && out2.valid) || (out8.to != out2.to)) && (!(out8.valid && out3.valid) || (out8.to != out3.to)) && (!(out8.valid && out4.valid) || (out8.to != out4.to)) && (!(out8.valid && out5.valid) || (out8.to != out5.to)) && (!(out8.valid && out6.valid) || (out8.to != out6.to)) && (!(out8.valid && out7.valid) || (out8.to != out7.to))
        && (!(out8.valid && out9.valid) || (out8.to != out9.to)) && (!(out8.valid && out10.valid) || (out8.to != out10.to)) && (!(out8.valid && out11.valid) || (out8.to != out11.to)) && (!(out8.valid && out12.valid) || (out8.to != out12.to)) && (!(out8.valid && out13.valid) || (out8.to != out13.to)) && (!(out8.valid && out14.valid) || (out8.to != out14.to)) && (!(out8.valid && out15.valid) || (out8.to != out15.to)) && (!(out9.valid && out0.valid) || (out9.to != out0.to)) && (!(out9.valid && out1.valid) || (out9.to != out1.to)) && (!(out9.valid && out2.valid) || (out9.to != out2.to)) && (!(out9.valid && out3.valid) || (out9.to != out3.to)) && (!(out9.valid && out4.valid) || (out9.to != out4.to)) && (!(out9.valid && out5.valid) || (out9.to != out5.to)) && (!(out9.valid && out6.valid) || (out9.to != out6.to)) && (!(out9.valid && out7.valid) || (out9.to != out7.to)) && (!(out9.valid && out8.valid) || (out9.to != out8.to)) && (!(out9.valid && out10.valid) || (out9.to != out10.to)) && (!(out9.valid && out11.valid) || (out9.to != out11.to)) && (!(out9.valid && out12.valid) || (out9.to != out12.to)) && (!(out9.valid && out13.valid) || (out9.to != out13.to)) && (!(out9.valid && out14.valid) || (out9.to != out14.to)) && (!(out9.valid && out15.valid) || (out9.to != out15.to)) && (!(out10.valid && out0.valid) || (out10.to != out0.to)) && (!(out10.valid && out1.valid) || (out10.to != out1.to)) && (!(out10.valid && out2.valid) || (out10.to != out2.to)) && (!(out10.valid && out3.valid) || (out10.to != out3.to)) && (!(out10.valid && out4.valid) || (out10.to != out4.to)) && (!(out10.valid && out5.valid) || (out10.to != out5.to)) && (!(out10.valid && out6.valid) || (out10.to != out6.to)) && (!(out10.valid && out7.valid) || (out10.to != out7.to)) && (!(out10.valid && out8.valid) || (out10.to != out8.to)) && (!(out10.valid && out9.valid) || (out10.to != out9.to)) && (!(out10.valid && out11.valid) || (out10.to != out11.to)) && (!(out10.valid && out12.valid) || (out10.to != out12.to)) && (!(out10.valid && out13.valid) || (out10.to != out13.to)) && (!(out10.valid && out14.valid) || (out10.to != out14.to)) && (!(out10.valid && out15.valid) || (out10.to != out15.to)) && (!(out11.valid && out0.valid) || (out11.to != out0.to)) && (!(out11.valid && out1.valid) || (out11.to != out1.to)) && (!(out11.valid && out2.valid) || (out11.to != out2.to)) && (!(out11.valid && out3.valid) || (out11.to != out3.to)) && (!(out11.valid && out4.valid) || (out11.to != out4.to)) && (!(out11.valid && out5.valid) || (out11.to != out5.to)) && (!(out11.valid && out6.valid) || (out11.to != out6.to)) && (!(out11.valid && out7.valid) || (out11.to != out7.to)) && (!(out11.valid && out8.valid) || (out11.to != out8.to)) && (!(out11.valid && out9.valid) || (out11.to != out9.to)) && (!(out11.valid && out10.valid) || (out11.to != out10.to)) && (!(out11.valid && out12.valid) || (out11.to != out12.to)) && (!(out11.valid && out13.valid) || (out11.to != out13.to)) && (!(out11.valid && out14.valid) || (out11.to != out14.to)) && (!(out11.valid && out15.valid) || (out11.to != out15.to)) && (!(out12.valid && out0.valid) || (out12.to != out0.to)) && (!(out12.valid && out1.valid) || (out12.to != out1.to)) && (!(out12.valid && out2.valid) || (out12.to != out2.to)) && (!(out12.valid && out3.valid) || (out12.to != out3.to)) && (!(out12.valid && out4.valid) || (out12.to != out4.to)) && (!(out12.valid && out5.valid) || (out12.to != out5.to)) && (!(out12.valid && out6.valid) || (out12.to != out6.to)) && (!(out12.valid && out7.valid) || (out12.to != out7.to)) && (!(out12.valid && out8.valid) || (out12.to != out8.to)) && (!(out12.valid && out9.valid) || (out12.to != out9.to)) && (!(out12.valid && out10.valid) || (out12.to != out10.to)) && (!(out12.valid && out11.valid) || (out12.to != out11.to)) && (!(out12.valid && out13.valid) || (out12.to != out13.to)) && (!(out12.valid && out14.valid) || (out12.to != out14.to)) && (!(out12.valid && out15.valid) || (out12.to != out15.to)) && (!(out13.valid && out0.valid) || (out13.to != out0.to)) && (!(out13.valid && out1.valid) || (out13.to != out1.to)) && (!(out13.valid && out2.valid) || (out13.to != out2.to)) && (!(out13.valid && out3.valid) || (out13.to != out3.to)) && (!(out13.valid && out4.valid) || (out13.to != out4.to)) && (!(out13.valid && out5.valid) || (out13.to != out5.to)) && (!(out13.valid && out6.valid) || (out13.to != out6.to)) && (!(out13.valid && out7.valid) || (out13.to != out7.to)) && (!(out13.valid && out8.valid) || (out13.to != out8.to)) && (!(out13.valid && out9.valid) || (out13.to != out9.to)) && (!(out13.valid && out10.valid) || (out13.to != out10.to)) && (!(out13.valid && out11.valid) || (out13.to != out11.to)) && (!(out13.valid && out12.valid) || (out13.to != out12.to)) && (!(out13.valid && out14.valid) || (out13.to != out14.to)) && (!(out13.valid && out15.valid) || (out13.to != out15.to)) && (!(out14.valid && out0.valid) || (out14.to != out0.to)) && (!(out14.valid && out1.valid) || (out14.to != out1.to)) && (!(out14.valid && out2.valid) || (out14.to != out2.to)) && (!(out14.valid && out3.valid) || (out14.to != out3.to)) && (!(out14.valid && out4.valid) || (out14.to != out4.to)) && (!(out14.valid && out5.valid) || (out14.to != out5.to)) && (!(out14.valid && out6.valid) || (out14.to != out6.to)) && (!(out14.valid && out7.valid) || (out14.to != out7.to)) && (!(out14.valid && out8.valid) || (out14.to != out8.to)) && (!(out14.valid && out9.valid) || (out14.to != out9.to)) && (!(out14.valid && out10.valid) || (out14.to != out10.to)) && (!(out14.valid && out11.valid) || (out14.to != out11.to)) && (!(out14.valid && out12.valid) || (out14.to != out12.to)) && (!(out14.valid && out13.valid) || (out14.to != out13.to)) && (!(out14.valid && out15.valid) || (out14.to != out15.to)) && (!(out15.valid && out0.valid) || (out15.to != out0.to)) && (!(out15.valid && out1.valid) || (out15.to != out1.to)) && (!(out15.valid && out2.valid) || (out15.to != out2.to)) && (!(out15.valid && out3.valid) || (out15.to != out3.to)) && (!(out15.valid && out4.valid) || (out15.to != out4.to)) && (!(out15.valid && out5.valid) || (out15.to != out5.to)) && (!(out15.valid && out6.valid) || (out15.to != out6.to)) && (!(out15.valid && out7.valid) || (out15.to != out7.to)) && (!(out15.valid && out8.valid) || (out15.to != out8.to)) && (!(out15.valid && out9.valid) || (out15.to != out9.to)) && (!(out15.valid && out10.valid) || (out15.to != out10.to)) && (!(out15.valid && out11.valid) || (out15.to != out11.to)) && (!(out15.valid && out12.valid) || (out15.to != out12.to)) && (!(out15.valid && out13.valid) || (out15.to != out13.to)) && (!(out15.valid && out14.valid) || (out15.to != out14.to)));
  correct_passthrough: assert property ((!out0.valid || ((in0.to == out0.to) && (in0.from == out0.from) &&
                         (in0.valid == out0.valid) && (in0.data == out0.data))) && (!out1.valid || ((in1.to == out1.to) && (in1.from == out1.from) &&
                         (in1.valid == out1.valid) && (in1.data == out1.data))) && (!out2.valid || ((in2.to == out2.to) && (in2.from == out2.from) &&
                         (in2.valid == out2.valid) && (in2.data == out2.data))) && (!out3.valid || ((in3.to == out3.to) && (in3.from == out3.from) &&
                         (in3.valid == out3.valid) && (in3.data == out3.data))) && (!out4.valid || ((in4.to == out4.to) && (in4.from == out4.from) &&
                         (in4.valid == out4.valid) && (in4.data == out4.data))) && (!out5.valid || ((in5.to == out5.to) && (in5.from == out5.from) &&
                         (in5.valid == out5.valid) && (in5.data == out5.data))) && (!out6.valid || ((in6.to == out6.to) && (in6.from == out6.from) &&
                         (in6.valid == out6.valid) && (in6.data == out6.data))) && (!out7.valid || ((in7.to == out7.to) && (in7.from == out7.from) &&
                         (in7.valid == out7.valid) && (in7.data == out7.data))) && (!out8.valid || ((in8.to == out8.to) && (in8.from == out8.from) &&
                         (in8.valid == out8.valid) && (in8.data == out8.data))) && (!out9.valid || ((in9.to == out9.to) && (in9.from == out9.from) &&
                         (in9.valid == out9.valid) && (in9.data == out9.data))) && (!out10.valid || ((in10.to == out10.to) && (in10.from == out10.from) &&
                         (in10.valid == out10.valid) && (in10.data == out10.data))) && (!out11.valid || ((in11.to == out11.to) && (in11.from == out11.from) &&
                         (in11.valid == out11.valid) && (in11.data == out11.data))) && (!out12.valid || ((in12.to == out12.to) && (in12.from == out12.from) &&
                         (in12.valid == out12.valid) && (in12.data == out12.data))) && (!out13.valid || ((in13.to == out13.to) && (in13.from == out13.from) &&
                         (in13.valid == out13.valid) && (in13.data == out13.data))) && (!out14.valid || ((in14.to == out14.to) && (in14.from == out14.from) &&
                         (in14.valid == out14.valid) && (in14.data == out14.data))) && (!out15.valid || ((in15.to == out15.to) && (in15.from == out15.from) &&
                         (in15.valid == out15.valid) && (in15.data == out15.data))));
  ack_when_forwareded: assert property ((!out0.valid || in0.ack) && (!out1.valid || in1.ack) && (!out2.valid || in2.ack) && (!out3.valid || in3.ack) && (!out4.valid || in4.ack) && (!out5.valid || in5.ack) && (!out6.valid || in6.ack) && (!out7.valid || in7.ack) && (!out8.valid || in8.ack) && (!out9.valid || in9.ack) && (!out10.valid || in10.ack) && (!out11.valid || in11.ack) && (!out12.valid || in12.ack) && (!out13.valid || in13.ack) && (!out14.valid || in14.ack) && (!out15.valid || in15.ack));
`endif
endmodule
