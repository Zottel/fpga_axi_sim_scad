`default_nettype none

module mib_simple_output_demux_14 (input wire [4-1:0] move_buffer_addr, input wire [4-1:0] immediate_buffer_addr, instruction_input_interface.consumer input_instr, instruction_input_interface.producer input_buffer_0, instruction_input_interface.producer input_buffer_1, instruction_input_interface.producer input_buffer_2, instruction_input_interface.producer input_buffer_3, instruction_input_interface.producer input_buffer_4, instruction_input_interface.producer input_buffer_5, instruction_input_interface.producer input_buffer_6, instruction_input_interface.producer input_buffer_7, instruction_input_interface.producer input_buffer_8, instruction_input_interface.producer input_buffer_9, instruction_input_interface.producer input_buffer_10, instruction_input_interface.producer input_buffer_11, instruction_input_interface.producer input_buffer_12, instruction_input_interface.producer input_buffer_13);
  assign input_buffer_0.move_from = (move_buffer_addr == 4'd0) ? input_instr.move_from : 0;
  assign input_buffer_0.move_valid = (move_buffer_addr == 4'd0) ? input_instr.move_valid : 0;
  assign input_buffer_1.move_from = (move_buffer_addr == 4'd1) ? input_instr.move_from : 0;
  assign input_buffer_1.move_valid = (move_buffer_addr == 4'd1) ? input_instr.move_valid : 0;
  assign input_buffer_2.move_from = (move_buffer_addr == 4'd2) ? input_instr.move_from : 0;
  assign input_buffer_2.move_valid = (move_buffer_addr == 4'd2) ? input_instr.move_valid : 0;
  assign input_buffer_3.move_from = (move_buffer_addr == 4'd3) ? input_instr.move_from : 0;
  assign input_buffer_3.move_valid = (move_buffer_addr == 4'd3) ? input_instr.move_valid : 0;
  assign input_buffer_4.move_from = (move_buffer_addr == 4'd4) ? input_instr.move_from : 0;
  assign input_buffer_4.move_valid = (move_buffer_addr == 4'd4) ? input_instr.move_valid : 0;
  assign input_buffer_5.move_from = (move_buffer_addr == 4'd5) ? input_instr.move_from : 0;
  assign input_buffer_5.move_valid = (move_buffer_addr == 4'd5) ? input_instr.move_valid : 0;
  assign input_buffer_6.move_from = (move_buffer_addr == 4'd6) ? input_instr.move_from : 0;
  assign input_buffer_6.move_valid = (move_buffer_addr == 4'd6) ? input_instr.move_valid : 0;
  assign input_buffer_7.move_from = (move_buffer_addr == 4'd7) ? input_instr.move_from : 0;
  assign input_buffer_7.move_valid = (move_buffer_addr == 4'd7) ? input_instr.move_valid : 0;
  assign input_buffer_8.move_from = (move_buffer_addr == 4'd8) ? input_instr.move_from : 0;
  assign input_buffer_8.move_valid = (move_buffer_addr == 4'd8) ? input_instr.move_valid : 0;
  assign input_buffer_9.move_from = (move_buffer_addr == 4'd9) ? input_instr.move_from : 0;
  assign input_buffer_9.move_valid = (move_buffer_addr == 4'd9) ? input_instr.move_valid : 0;
  assign input_buffer_10.move_from = (move_buffer_addr == 4'd10) ? input_instr.move_from : 0;
  assign input_buffer_10.move_valid = (move_buffer_addr == 4'd10) ? input_instr.move_valid : 0;
  assign input_buffer_11.move_from = (move_buffer_addr == 4'd11) ? input_instr.move_from : 0;
  assign input_buffer_11.move_valid = (move_buffer_addr == 4'd11) ? input_instr.move_valid : 0;
  assign input_buffer_12.move_from = (move_buffer_addr == 4'd12) ? input_instr.move_from : 0;
  assign input_buffer_12.move_valid = (move_buffer_addr == 4'd12) ? input_instr.move_valid : 0;
  assign input_buffer_13.move_from = (move_buffer_addr == 4'd13) ? input_instr.move_from : 0;
  assign input_buffer_13.move_valid = (move_buffer_addr == 4'd13) ? input_instr.move_valid : 0;
assign input_instr.move_ack = (move_buffer_addr == {4{1'b1}})||((move_buffer_addr == 4'd0) && input_buffer_0.move_ack)||((move_buffer_addr == 4'd1) && input_buffer_1.move_ack)||((move_buffer_addr == 4'd2) && input_buffer_2.move_ack)||((move_buffer_addr == 4'd3) && input_buffer_3.move_ack)||((move_buffer_addr == 4'd4) && input_buffer_4.move_ack)||((move_buffer_addr == 4'd5) && input_buffer_5.move_ack)||((move_buffer_addr == 4'd6) && input_buffer_6.move_ack)||((move_buffer_addr == 4'd7) && input_buffer_7.move_ack)||((move_buffer_addr == 4'd8) && input_buffer_8.move_ack)||((move_buffer_addr == 4'd9) && input_buffer_9.move_ack)||((move_buffer_addr == 4'd10) && input_buffer_10.move_ack)||((move_buffer_addr == 4'd11) && input_buffer_11.move_ack)||((move_buffer_addr == 4'd12) && input_buffer_12.move_ack)||((move_buffer_addr == 4'd13) && input_buffer_13.move_ack);
  assign input_buffer_0.immediate = (immediate_buffer_addr == 4'd0) ? input_instr.immediate : 0;
  assign input_buffer_0.immediate_valid = (immediate_buffer_addr == 4'd0) ? input_instr.immediate_valid : 0;
  assign input_buffer_1.immediate = (immediate_buffer_addr == 4'd1) ? input_instr.immediate : 0;
  assign input_buffer_1.immediate_valid = (immediate_buffer_addr == 4'd1) ? input_instr.immediate_valid : 0;
  assign input_buffer_2.immediate = (immediate_buffer_addr == 4'd2) ? input_instr.immediate : 0;
  assign input_buffer_2.immediate_valid = (immediate_buffer_addr == 4'd2) ? input_instr.immediate_valid : 0;
  assign input_buffer_3.immediate = (immediate_buffer_addr == 4'd3) ? input_instr.immediate : 0;
  assign input_buffer_3.immediate_valid = (immediate_buffer_addr == 4'd3) ? input_instr.immediate_valid : 0;
  assign input_buffer_4.immediate = (immediate_buffer_addr == 4'd4) ? input_instr.immediate : 0;
  assign input_buffer_4.immediate_valid = (immediate_buffer_addr == 4'd4) ? input_instr.immediate_valid : 0;
  assign input_buffer_5.immediate = (immediate_buffer_addr == 4'd5) ? input_instr.immediate : 0;
  assign input_buffer_5.immediate_valid = (immediate_buffer_addr == 4'd5) ? input_instr.immediate_valid : 0;
  assign input_buffer_6.immediate = (immediate_buffer_addr == 4'd6) ? input_instr.immediate : 0;
  assign input_buffer_6.immediate_valid = (immediate_buffer_addr == 4'd6) ? input_instr.immediate_valid : 0;
  assign input_buffer_7.immediate = (immediate_buffer_addr == 4'd7) ? input_instr.immediate : 0;
  assign input_buffer_7.immediate_valid = (immediate_buffer_addr == 4'd7) ? input_instr.immediate_valid : 0;
  assign input_buffer_8.immediate = (immediate_buffer_addr == 4'd8) ? input_instr.immediate : 0;
  assign input_buffer_8.immediate_valid = (immediate_buffer_addr == 4'd8) ? input_instr.immediate_valid : 0;
  assign input_buffer_9.immediate = (immediate_buffer_addr == 4'd9) ? input_instr.immediate : 0;
  assign input_buffer_9.immediate_valid = (immediate_buffer_addr == 4'd9) ? input_instr.immediate_valid : 0;
  assign input_buffer_10.immediate = (immediate_buffer_addr == 4'd10) ? input_instr.immediate : 0;
  assign input_buffer_10.immediate_valid = (immediate_buffer_addr == 4'd10) ? input_instr.immediate_valid : 0;
  assign input_buffer_11.immediate = (immediate_buffer_addr == 4'd11) ? input_instr.immediate : 0;
  assign input_buffer_11.immediate_valid = (immediate_buffer_addr == 4'd11) ? input_instr.immediate_valid : 0;
  assign input_buffer_12.immediate = (immediate_buffer_addr == 4'd12) ? input_instr.immediate : 0;
  assign input_buffer_12.immediate_valid = (immediate_buffer_addr == 4'd12) ? input_instr.immediate_valid : 0;
  assign input_buffer_13.immediate = (immediate_buffer_addr == 4'd13) ? input_instr.immediate : 0;
  assign input_buffer_13.immediate_valid = (immediate_buffer_addr == 4'd13) ? input_instr.immediate_valid : 0;
assign input_instr.immediate_ack = ((immediate_buffer_addr == 4'd0) && input_buffer_0.move_ack)||((immediate_buffer_addr == 4'd1) && input_buffer_1.move_ack)||((immediate_buffer_addr == 4'd2) && input_buffer_2.move_ack)||((immediate_buffer_addr == 4'd3) && input_buffer_3.move_ack)||((immediate_buffer_addr == 4'd4) && input_buffer_4.move_ack)||((immediate_buffer_addr == 4'd5) && input_buffer_5.move_ack)||((immediate_buffer_addr == 4'd6) && input_buffer_6.move_ack)||((immediate_buffer_addr == 4'd7) && input_buffer_7.move_ack)||((immediate_buffer_addr == 4'd8) && input_buffer_8.move_ack)||((immediate_buffer_addr == 4'd9) && input_buffer_9.move_ack)||((immediate_buffer_addr == 4'd10) && input_buffer_10.move_ack)||((immediate_buffer_addr == 4'd11) && input_buffer_11.move_ack)||((immediate_buffer_addr == 4'd12) && input_buffer_12.move_ack)||((immediate_buffer_addr == 4'd13) && input_buffer_13.move_ack);
endmodule
