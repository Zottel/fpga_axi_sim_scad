`default_nettype none

module TNT_BIN_HC0_JaSJ17_68_16_3 (
output wire [70-1:0] out0,
output wire [70-1:0] out1,
output wire [70-1:0] out2,
output wire [70-1:0] out3,
output wire [70-1:0] out4,
output wire [70-1:0] out5,
output wire [70-1:0] out6,
output wire [70-1:0] out7,
output wire [70-1:0] out8,
output wire [70-1:0] out9,
output wire [70-1:0] out10,
output wire [70-1:0] out11,
output wire [70-1:0] out12,
output wire [70-1:0] out13,
output wire [70-1:0] out14,
output wire [70-1:0] out15,
input wire [71-1:0] in0,
input wire [71-1:0] in1,
input wire [71-1:0] in2,
input wire [71-1:0] in3,
input wire [71-1:0] in4,
input wire [71-1:0] in5,
input wire [71-1:0] in6,
input wire [71-1:0] in7,
input wire [71-1:0] in8,
input wire [71-1:0] in9,
input wire [71-1:0] in10,
input wire [71-1:0] in11,
input wire [71-1:0] in12,
input wire [71-1:0] in13,
input wire [71-1:0] in14,
input wire [71-1:0] in15);
    wire x0_0;
    wire x0_1;
    wire x0_2;
    wire x0_3;
    wire x0_4;
    wire x0_5;
    wire x0_6;
    wire x0_7;
    wire x0_8;
    wire x0_9;
    wire x0_10;
    wire x0_11;
    wire x0_12;
    wire x0_13;
    wire x0_14;
    wire x0_15;
    wire x0_16;
    wire x0_17;
    wire x0_18;
    wire x0_19;
    wire x0_20;
    wire x0_21;
    wire x0_22;
    wire x0_23;
    wire x0_24;
    wire x0_25;
    wire x0_26;
    wire x0_27;
    wire x0_28;
    wire x0_29;
    wire x0_30;
    wire x0_31;
    wire x0_32;
    wire x0_33;
    wire x0_34;
    wire x0_35;
    wire x0_36;
    wire x0_37;
    wire x0_38;
    wire x0_39;
    wire x0_40;
    wire x0_41;
    wire x0_42;
    wire x0_43;
    wire x0_44;
    wire x0_45;
    wire x0_46;
    wire x0_47;
    wire x0_48;
    wire x0_49;
    wire x0_50;
    wire x0_51;
    wire x0_52;
    wire x0_53;
    wire x0_54;
    wire x0_55;
    wire x0_56;
    wire x0_57;
    wire x0_58;
    wire x0_59;
    wire x0_60;
    wire x0_61;
    wire x0_62;
    wire x0_63;
    wire x0_64;
    wire x0_65;
    wire x0_66;
    wire x0_67;
    wire x0_68;
    wire x0_69;
    wire x0_70;
    assign x0_0 = in0[0];
    assign x0_1 = in0[1];
    assign x0_2 = in0[2];
    assign x0_3 = in0[3];
    assign x0_4 = in0[4];
    assign x0_5 = in0[5];
    assign x0_6 = in0[6];
    assign x0_7 = in0[7];
    assign x0_8 = in0[8];
    assign x0_9 = in0[9];
    assign x0_10 = in0[10];
    assign x0_11 = in0[11];
    assign x0_12 = in0[12];
    assign x0_13 = in0[13];
    assign x0_14 = in0[14];
    assign x0_15 = in0[15];
    assign x0_16 = in0[16];
    assign x0_17 = in0[17];
    assign x0_18 = in0[18];
    assign x0_19 = in0[19];
    assign x0_20 = in0[20];
    assign x0_21 = in0[21];
    assign x0_22 = in0[22];
    assign x0_23 = in0[23];
    assign x0_24 = in0[24];
    assign x0_25 = in0[25];
    assign x0_26 = in0[26];
    assign x0_27 = in0[27];
    assign x0_28 = in0[28];
    assign x0_29 = in0[29];
    assign x0_30 = in0[30];
    assign x0_31 = in0[31];
    assign x0_32 = in0[32];
    assign x0_33 = in0[33];
    assign x0_34 = in0[34];
    assign x0_35 = in0[35];
    assign x0_36 = in0[36];
    assign x0_37 = in0[37];
    assign x0_38 = in0[38];
    assign x0_39 = in0[39];
    assign x0_40 = in0[40];
    assign x0_41 = in0[41];
    assign x0_42 = in0[42];
    assign x0_43 = in0[43];
    assign x0_44 = in0[44];
    assign x0_45 = in0[45];
    assign x0_46 = in0[46];
    assign x0_47 = in0[47];
    assign x0_48 = in0[48];
    assign x0_49 = in0[49];
    assign x0_50 = in0[50];
    assign x0_51 = in0[51];
    assign x0_52 = in0[52];
    assign x0_53 = in0[53];
    assign x0_54 = in0[54];
    assign x0_55 = in0[55];
    assign x0_56 = in0[56];
    assign x0_57 = in0[57];
    assign x0_58 = in0[58];
    assign x0_59 = in0[59];
    assign x0_60 = in0[60];
    assign x0_61 = in0[61];
    assign x0_62 = in0[62];
    assign x0_63 = in0[63];
    assign x0_64 = in0[64];
    assign x0_65 = in0[65];
    assign x0_66 = in0[66];
    assign x0_67 = in0[67];
    assign x0_68 = in0[68];
    assign x0_69 = in0[69];
    assign x0_70 = in0[70];
    wire x1_0;
    wire x1_1;
    wire x1_2;
    wire x1_3;
    wire x1_4;
    wire x1_5;
    wire x1_6;
    wire x1_7;
    wire x1_8;
    wire x1_9;
    wire x1_10;
    wire x1_11;
    wire x1_12;
    wire x1_13;
    wire x1_14;
    wire x1_15;
    wire x1_16;
    wire x1_17;
    wire x1_18;
    wire x1_19;
    wire x1_20;
    wire x1_21;
    wire x1_22;
    wire x1_23;
    wire x1_24;
    wire x1_25;
    wire x1_26;
    wire x1_27;
    wire x1_28;
    wire x1_29;
    wire x1_30;
    wire x1_31;
    wire x1_32;
    wire x1_33;
    wire x1_34;
    wire x1_35;
    wire x1_36;
    wire x1_37;
    wire x1_38;
    wire x1_39;
    wire x1_40;
    wire x1_41;
    wire x1_42;
    wire x1_43;
    wire x1_44;
    wire x1_45;
    wire x1_46;
    wire x1_47;
    wire x1_48;
    wire x1_49;
    wire x1_50;
    wire x1_51;
    wire x1_52;
    wire x1_53;
    wire x1_54;
    wire x1_55;
    wire x1_56;
    wire x1_57;
    wire x1_58;
    wire x1_59;
    wire x1_60;
    wire x1_61;
    wire x1_62;
    wire x1_63;
    wire x1_64;
    wire x1_65;
    wire x1_66;
    wire x1_67;
    wire x1_68;
    wire x1_69;
    wire x1_70;
    assign x1_0 = in1[0];
    assign x1_1 = in1[1];
    assign x1_2 = in1[2];
    assign x1_3 = in1[3];
    assign x1_4 = in1[4];
    assign x1_5 = in1[5];
    assign x1_6 = in1[6];
    assign x1_7 = in1[7];
    assign x1_8 = in1[8];
    assign x1_9 = in1[9];
    assign x1_10 = in1[10];
    assign x1_11 = in1[11];
    assign x1_12 = in1[12];
    assign x1_13 = in1[13];
    assign x1_14 = in1[14];
    assign x1_15 = in1[15];
    assign x1_16 = in1[16];
    assign x1_17 = in1[17];
    assign x1_18 = in1[18];
    assign x1_19 = in1[19];
    assign x1_20 = in1[20];
    assign x1_21 = in1[21];
    assign x1_22 = in1[22];
    assign x1_23 = in1[23];
    assign x1_24 = in1[24];
    assign x1_25 = in1[25];
    assign x1_26 = in1[26];
    assign x1_27 = in1[27];
    assign x1_28 = in1[28];
    assign x1_29 = in1[29];
    assign x1_30 = in1[30];
    assign x1_31 = in1[31];
    assign x1_32 = in1[32];
    assign x1_33 = in1[33];
    assign x1_34 = in1[34];
    assign x1_35 = in1[35];
    assign x1_36 = in1[36];
    assign x1_37 = in1[37];
    assign x1_38 = in1[38];
    assign x1_39 = in1[39];
    assign x1_40 = in1[40];
    assign x1_41 = in1[41];
    assign x1_42 = in1[42];
    assign x1_43 = in1[43];
    assign x1_44 = in1[44];
    assign x1_45 = in1[45];
    assign x1_46 = in1[46];
    assign x1_47 = in1[47];
    assign x1_48 = in1[48];
    assign x1_49 = in1[49];
    assign x1_50 = in1[50];
    assign x1_51 = in1[51];
    assign x1_52 = in1[52];
    assign x1_53 = in1[53];
    assign x1_54 = in1[54];
    assign x1_55 = in1[55];
    assign x1_56 = in1[56];
    assign x1_57 = in1[57];
    assign x1_58 = in1[58];
    assign x1_59 = in1[59];
    assign x1_60 = in1[60];
    assign x1_61 = in1[61];
    assign x1_62 = in1[62];
    assign x1_63 = in1[63];
    assign x1_64 = in1[64];
    assign x1_65 = in1[65];
    assign x1_66 = in1[66];
    assign x1_67 = in1[67];
    assign x1_68 = in1[68];
    assign x1_69 = in1[69];
    assign x1_70 = in1[70];
    wire x2_0;
    wire x2_1;
    wire x2_2;
    wire x2_3;
    wire x2_4;
    wire x2_5;
    wire x2_6;
    wire x2_7;
    wire x2_8;
    wire x2_9;
    wire x2_10;
    wire x2_11;
    wire x2_12;
    wire x2_13;
    wire x2_14;
    wire x2_15;
    wire x2_16;
    wire x2_17;
    wire x2_18;
    wire x2_19;
    wire x2_20;
    wire x2_21;
    wire x2_22;
    wire x2_23;
    wire x2_24;
    wire x2_25;
    wire x2_26;
    wire x2_27;
    wire x2_28;
    wire x2_29;
    wire x2_30;
    wire x2_31;
    wire x2_32;
    wire x2_33;
    wire x2_34;
    wire x2_35;
    wire x2_36;
    wire x2_37;
    wire x2_38;
    wire x2_39;
    wire x2_40;
    wire x2_41;
    wire x2_42;
    wire x2_43;
    wire x2_44;
    wire x2_45;
    wire x2_46;
    wire x2_47;
    wire x2_48;
    wire x2_49;
    wire x2_50;
    wire x2_51;
    wire x2_52;
    wire x2_53;
    wire x2_54;
    wire x2_55;
    wire x2_56;
    wire x2_57;
    wire x2_58;
    wire x2_59;
    wire x2_60;
    wire x2_61;
    wire x2_62;
    wire x2_63;
    wire x2_64;
    wire x2_65;
    wire x2_66;
    wire x2_67;
    wire x2_68;
    wire x2_69;
    wire x2_70;
    assign x2_0 = in2[0];
    assign x2_1 = in2[1];
    assign x2_2 = in2[2];
    assign x2_3 = in2[3];
    assign x2_4 = in2[4];
    assign x2_5 = in2[5];
    assign x2_6 = in2[6];
    assign x2_7 = in2[7];
    assign x2_8 = in2[8];
    assign x2_9 = in2[9];
    assign x2_10 = in2[10];
    assign x2_11 = in2[11];
    assign x2_12 = in2[12];
    assign x2_13 = in2[13];
    assign x2_14 = in2[14];
    assign x2_15 = in2[15];
    assign x2_16 = in2[16];
    assign x2_17 = in2[17];
    assign x2_18 = in2[18];
    assign x2_19 = in2[19];
    assign x2_20 = in2[20];
    assign x2_21 = in2[21];
    assign x2_22 = in2[22];
    assign x2_23 = in2[23];
    assign x2_24 = in2[24];
    assign x2_25 = in2[25];
    assign x2_26 = in2[26];
    assign x2_27 = in2[27];
    assign x2_28 = in2[28];
    assign x2_29 = in2[29];
    assign x2_30 = in2[30];
    assign x2_31 = in2[31];
    assign x2_32 = in2[32];
    assign x2_33 = in2[33];
    assign x2_34 = in2[34];
    assign x2_35 = in2[35];
    assign x2_36 = in2[36];
    assign x2_37 = in2[37];
    assign x2_38 = in2[38];
    assign x2_39 = in2[39];
    assign x2_40 = in2[40];
    assign x2_41 = in2[41];
    assign x2_42 = in2[42];
    assign x2_43 = in2[43];
    assign x2_44 = in2[44];
    assign x2_45 = in2[45];
    assign x2_46 = in2[46];
    assign x2_47 = in2[47];
    assign x2_48 = in2[48];
    assign x2_49 = in2[49];
    assign x2_50 = in2[50];
    assign x2_51 = in2[51];
    assign x2_52 = in2[52];
    assign x2_53 = in2[53];
    assign x2_54 = in2[54];
    assign x2_55 = in2[55];
    assign x2_56 = in2[56];
    assign x2_57 = in2[57];
    assign x2_58 = in2[58];
    assign x2_59 = in2[59];
    assign x2_60 = in2[60];
    assign x2_61 = in2[61];
    assign x2_62 = in2[62];
    assign x2_63 = in2[63];
    assign x2_64 = in2[64];
    assign x2_65 = in2[65];
    assign x2_66 = in2[66];
    assign x2_67 = in2[67];
    assign x2_68 = in2[68];
    assign x2_69 = in2[69];
    assign x2_70 = in2[70];
    wire x3_0;
    wire x3_1;
    wire x3_2;
    wire x3_3;
    wire x3_4;
    wire x3_5;
    wire x3_6;
    wire x3_7;
    wire x3_8;
    wire x3_9;
    wire x3_10;
    wire x3_11;
    wire x3_12;
    wire x3_13;
    wire x3_14;
    wire x3_15;
    wire x3_16;
    wire x3_17;
    wire x3_18;
    wire x3_19;
    wire x3_20;
    wire x3_21;
    wire x3_22;
    wire x3_23;
    wire x3_24;
    wire x3_25;
    wire x3_26;
    wire x3_27;
    wire x3_28;
    wire x3_29;
    wire x3_30;
    wire x3_31;
    wire x3_32;
    wire x3_33;
    wire x3_34;
    wire x3_35;
    wire x3_36;
    wire x3_37;
    wire x3_38;
    wire x3_39;
    wire x3_40;
    wire x3_41;
    wire x3_42;
    wire x3_43;
    wire x3_44;
    wire x3_45;
    wire x3_46;
    wire x3_47;
    wire x3_48;
    wire x3_49;
    wire x3_50;
    wire x3_51;
    wire x3_52;
    wire x3_53;
    wire x3_54;
    wire x3_55;
    wire x3_56;
    wire x3_57;
    wire x3_58;
    wire x3_59;
    wire x3_60;
    wire x3_61;
    wire x3_62;
    wire x3_63;
    wire x3_64;
    wire x3_65;
    wire x3_66;
    wire x3_67;
    wire x3_68;
    wire x3_69;
    wire x3_70;
    assign x3_0 = in3[0];
    assign x3_1 = in3[1];
    assign x3_2 = in3[2];
    assign x3_3 = in3[3];
    assign x3_4 = in3[4];
    assign x3_5 = in3[5];
    assign x3_6 = in3[6];
    assign x3_7 = in3[7];
    assign x3_8 = in3[8];
    assign x3_9 = in3[9];
    assign x3_10 = in3[10];
    assign x3_11 = in3[11];
    assign x3_12 = in3[12];
    assign x3_13 = in3[13];
    assign x3_14 = in3[14];
    assign x3_15 = in3[15];
    assign x3_16 = in3[16];
    assign x3_17 = in3[17];
    assign x3_18 = in3[18];
    assign x3_19 = in3[19];
    assign x3_20 = in3[20];
    assign x3_21 = in3[21];
    assign x3_22 = in3[22];
    assign x3_23 = in3[23];
    assign x3_24 = in3[24];
    assign x3_25 = in3[25];
    assign x3_26 = in3[26];
    assign x3_27 = in3[27];
    assign x3_28 = in3[28];
    assign x3_29 = in3[29];
    assign x3_30 = in3[30];
    assign x3_31 = in3[31];
    assign x3_32 = in3[32];
    assign x3_33 = in3[33];
    assign x3_34 = in3[34];
    assign x3_35 = in3[35];
    assign x3_36 = in3[36];
    assign x3_37 = in3[37];
    assign x3_38 = in3[38];
    assign x3_39 = in3[39];
    assign x3_40 = in3[40];
    assign x3_41 = in3[41];
    assign x3_42 = in3[42];
    assign x3_43 = in3[43];
    assign x3_44 = in3[44];
    assign x3_45 = in3[45];
    assign x3_46 = in3[46];
    assign x3_47 = in3[47];
    assign x3_48 = in3[48];
    assign x3_49 = in3[49];
    assign x3_50 = in3[50];
    assign x3_51 = in3[51];
    assign x3_52 = in3[52];
    assign x3_53 = in3[53];
    assign x3_54 = in3[54];
    assign x3_55 = in3[55];
    assign x3_56 = in3[56];
    assign x3_57 = in3[57];
    assign x3_58 = in3[58];
    assign x3_59 = in3[59];
    assign x3_60 = in3[60];
    assign x3_61 = in3[61];
    assign x3_62 = in3[62];
    assign x3_63 = in3[63];
    assign x3_64 = in3[64];
    assign x3_65 = in3[65];
    assign x3_66 = in3[66];
    assign x3_67 = in3[67];
    assign x3_68 = in3[68];
    assign x3_69 = in3[69];
    assign x3_70 = in3[70];
    wire x4_0;
    wire x4_1;
    wire x4_2;
    wire x4_3;
    wire x4_4;
    wire x4_5;
    wire x4_6;
    wire x4_7;
    wire x4_8;
    wire x4_9;
    wire x4_10;
    wire x4_11;
    wire x4_12;
    wire x4_13;
    wire x4_14;
    wire x4_15;
    wire x4_16;
    wire x4_17;
    wire x4_18;
    wire x4_19;
    wire x4_20;
    wire x4_21;
    wire x4_22;
    wire x4_23;
    wire x4_24;
    wire x4_25;
    wire x4_26;
    wire x4_27;
    wire x4_28;
    wire x4_29;
    wire x4_30;
    wire x4_31;
    wire x4_32;
    wire x4_33;
    wire x4_34;
    wire x4_35;
    wire x4_36;
    wire x4_37;
    wire x4_38;
    wire x4_39;
    wire x4_40;
    wire x4_41;
    wire x4_42;
    wire x4_43;
    wire x4_44;
    wire x4_45;
    wire x4_46;
    wire x4_47;
    wire x4_48;
    wire x4_49;
    wire x4_50;
    wire x4_51;
    wire x4_52;
    wire x4_53;
    wire x4_54;
    wire x4_55;
    wire x4_56;
    wire x4_57;
    wire x4_58;
    wire x4_59;
    wire x4_60;
    wire x4_61;
    wire x4_62;
    wire x4_63;
    wire x4_64;
    wire x4_65;
    wire x4_66;
    wire x4_67;
    wire x4_68;
    wire x4_69;
    wire x4_70;
    assign x4_0 = in4[0];
    assign x4_1 = in4[1];
    assign x4_2 = in4[2];
    assign x4_3 = in4[3];
    assign x4_4 = in4[4];
    assign x4_5 = in4[5];
    assign x4_6 = in4[6];
    assign x4_7 = in4[7];
    assign x4_8 = in4[8];
    assign x4_9 = in4[9];
    assign x4_10 = in4[10];
    assign x4_11 = in4[11];
    assign x4_12 = in4[12];
    assign x4_13 = in4[13];
    assign x4_14 = in4[14];
    assign x4_15 = in4[15];
    assign x4_16 = in4[16];
    assign x4_17 = in4[17];
    assign x4_18 = in4[18];
    assign x4_19 = in4[19];
    assign x4_20 = in4[20];
    assign x4_21 = in4[21];
    assign x4_22 = in4[22];
    assign x4_23 = in4[23];
    assign x4_24 = in4[24];
    assign x4_25 = in4[25];
    assign x4_26 = in4[26];
    assign x4_27 = in4[27];
    assign x4_28 = in4[28];
    assign x4_29 = in4[29];
    assign x4_30 = in4[30];
    assign x4_31 = in4[31];
    assign x4_32 = in4[32];
    assign x4_33 = in4[33];
    assign x4_34 = in4[34];
    assign x4_35 = in4[35];
    assign x4_36 = in4[36];
    assign x4_37 = in4[37];
    assign x4_38 = in4[38];
    assign x4_39 = in4[39];
    assign x4_40 = in4[40];
    assign x4_41 = in4[41];
    assign x4_42 = in4[42];
    assign x4_43 = in4[43];
    assign x4_44 = in4[44];
    assign x4_45 = in4[45];
    assign x4_46 = in4[46];
    assign x4_47 = in4[47];
    assign x4_48 = in4[48];
    assign x4_49 = in4[49];
    assign x4_50 = in4[50];
    assign x4_51 = in4[51];
    assign x4_52 = in4[52];
    assign x4_53 = in4[53];
    assign x4_54 = in4[54];
    assign x4_55 = in4[55];
    assign x4_56 = in4[56];
    assign x4_57 = in4[57];
    assign x4_58 = in4[58];
    assign x4_59 = in4[59];
    assign x4_60 = in4[60];
    assign x4_61 = in4[61];
    assign x4_62 = in4[62];
    assign x4_63 = in4[63];
    assign x4_64 = in4[64];
    assign x4_65 = in4[65];
    assign x4_66 = in4[66];
    assign x4_67 = in4[67];
    assign x4_68 = in4[68];
    assign x4_69 = in4[69];
    assign x4_70 = in4[70];
    wire x5_0;
    wire x5_1;
    wire x5_2;
    wire x5_3;
    wire x5_4;
    wire x5_5;
    wire x5_6;
    wire x5_7;
    wire x5_8;
    wire x5_9;
    wire x5_10;
    wire x5_11;
    wire x5_12;
    wire x5_13;
    wire x5_14;
    wire x5_15;
    wire x5_16;
    wire x5_17;
    wire x5_18;
    wire x5_19;
    wire x5_20;
    wire x5_21;
    wire x5_22;
    wire x5_23;
    wire x5_24;
    wire x5_25;
    wire x5_26;
    wire x5_27;
    wire x5_28;
    wire x5_29;
    wire x5_30;
    wire x5_31;
    wire x5_32;
    wire x5_33;
    wire x5_34;
    wire x5_35;
    wire x5_36;
    wire x5_37;
    wire x5_38;
    wire x5_39;
    wire x5_40;
    wire x5_41;
    wire x5_42;
    wire x5_43;
    wire x5_44;
    wire x5_45;
    wire x5_46;
    wire x5_47;
    wire x5_48;
    wire x5_49;
    wire x5_50;
    wire x5_51;
    wire x5_52;
    wire x5_53;
    wire x5_54;
    wire x5_55;
    wire x5_56;
    wire x5_57;
    wire x5_58;
    wire x5_59;
    wire x5_60;
    wire x5_61;
    wire x5_62;
    wire x5_63;
    wire x5_64;
    wire x5_65;
    wire x5_66;
    wire x5_67;
    wire x5_68;
    wire x5_69;
    wire x5_70;
    assign x5_0 = in5[0];
    assign x5_1 = in5[1];
    assign x5_2 = in5[2];
    assign x5_3 = in5[3];
    assign x5_4 = in5[4];
    assign x5_5 = in5[5];
    assign x5_6 = in5[6];
    assign x5_7 = in5[7];
    assign x5_8 = in5[8];
    assign x5_9 = in5[9];
    assign x5_10 = in5[10];
    assign x5_11 = in5[11];
    assign x5_12 = in5[12];
    assign x5_13 = in5[13];
    assign x5_14 = in5[14];
    assign x5_15 = in5[15];
    assign x5_16 = in5[16];
    assign x5_17 = in5[17];
    assign x5_18 = in5[18];
    assign x5_19 = in5[19];
    assign x5_20 = in5[20];
    assign x5_21 = in5[21];
    assign x5_22 = in5[22];
    assign x5_23 = in5[23];
    assign x5_24 = in5[24];
    assign x5_25 = in5[25];
    assign x5_26 = in5[26];
    assign x5_27 = in5[27];
    assign x5_28 = in5[28];
    assign x5_29 = in5[29];
    assign x5_30 = in5[30];
    assign x5_31 = in5[31];
    assign x5_32 = in5[32];
    assign x5_33 = in5[33];
    assign x5_34 = in5[34];
    assign x5_35 = in5[35];
    assign x5_36 = in5[36];
    assign x5_37 = in5[37];
    assign x5_38 = in5[38];
    assign x5_39 = in5[39];
    assign x5_40 = in5[40];
    assign x5_41 = in5[41];
    assign x5_42 = in5[42];
    assign x5_43 = in5[43];
    assign x5_44 = in5[44];
    assign x5_45 = in5[45];
    assign x5_46 = in5[46];
    assign x5_47 = in5[47];
    assign x5_48 = in5[48];
    assign x5_49 = in5[49];
    assign x5_50 = in5[50];
    assign x5_51 = in5[51];
    assign x5_52 = in5[52];
    assign x5_53 = in5[53];
    assign x5_54 = in5[54];
    assign x5_55 = in5[55];
    assign x5_56 = in5[56];
    assign x5_57 = in5[57];
    assign x5_58 = in5[58];
    assign x5_59 = in5[59];
    assign x5_60 = in5[60];
    assign x5_61 = in5[61];
    assign x5_62 = in5[62];
    assign x5_63 = in5[63];
    assign x5_64 = in5[64];
    assign x5_65 = in5[65];
    assign x5_66 = in5[66];
    assign x5_67 = in5[67];
    assign x5_68 = in5[68];
    assign x5_69 = in5[69];
    assign x5_70 = in5[70];
    wire x6_0;
    wire x6_1;
    wire x6_2;
    wire x6_3;
    wire x6_4;
    wire x6_5;
    wire x6_6;
    wire x6_7;
    wire x6_8;
    wire x6_9;
    wire x6_10;
    wire x6_11;
    wire x6_12;
    wire x6_13;
    wire x6_14;
    wire x6_15;
    wire x6_16;
    wire x6_17;
    wire x6_18;
    wire x6_19;
    wire x6_20;
    wire x6_21;
    wire x6_22;
    wire x6_23;
    wire x6_24;
    wire x6_25;
    wire x6_26;
    wire x6_27;
    wire x6_28;
    wire x6_29;
    wire x6_30;
    wire x6_31;
    wire x6_32;
    wire x6_33;
    wire x6_34;
    wire x6_35;
    wire x6_36;
    wire x6_37;
    wire x6_38;
    wire x6_39;
    wire x6_40;
    wire x6_41;
    wire x6_42;
    wire x6_43;
    wire x6_44;
    wire x6_45;
    wire x6_46;
    wire x6_47;
    wire x6_48;
    wire x6_49;
    wire x6_50;
    wire x6_51;
    wire x6_52;
    wire x6_53;
    wire x6_54;
    wire x6_55;
    wire x6_56;
    wire x6_57;
    wire x6_58;
    wire x6_59;
    wire x6_60;
    wire x6_61;
    wire x6_62;
    wire x6_63;
    wire x6_64;
    wire x6_65;
    wire x6_66;
    wire x6_67;
    wire x6_68;
    wire x6_69;
    wire x6_70;
    assign x6_0 = in6[0];
    assign x6_1 = in6[1];
    assign x6_2 = in6[2];
    assign x6_3 = in6[3];
    assign x6_4 = in6[4];
    assign x6_5 = in6[5];
    assign x6_6 = in6[6];
    assign x6_7 = in6[7];
    assign x6_8 = in6[8];
    assign x6_9 = in6[9];
    assign x6_10 = in6[10];
    assign x6_11 = in6[11];
    assign x6_12 = in6[12];
    assign x6_13 = in6[13];
    assign x6_14 = in6[14];
    assign x6_15 = in6[15];
    assign x6_16 = in6[16];
    assign x6_17 = in6[17];
    assign x6_18 = in6[18];
    assign x6_19 = in6[19];
    assign x6_20 = in6[20];
    assign x6_21 = in6[21];
    assign x6_22 = in6[22];
    assign x6_23 = in6[23];
    assign x6_24 = in6[24];
    assign x6_25 = in6[25];
    assign x6_26 = in6[26];
    assign x6_27 = in6[27];
    assign x6_28 = in6[28];
    assign x6_29 = in6[29];
    assign x6_30 = in6[30];
    assign x6_31 = in6[31];
    assign x6_32 = in6[32];
    assign x6_33 = in6[33];
    assign x6_34 = in6[34];
    assign x6_35 = in6[35];
    assign x6_36 = in6[36];
    assign x6_37 = in6[37];
    assign x6_38 = in6[38];
    assign x6_39 = in6[39];
    assign x6_40 = in6[40];
    assign x6_41 = in6[41];
    assign x6_42 = in6[42];
    assign x6_43 = in6[43];
    assign x6_44 = in6[44];
    assign x6_45 = in6[45];
    assign x6_46 = in6[46];
    assign x6_47 = in6[47];
    assign x6_48 = in6[48];
    assign x6_49 = in6[49];
    assign x6_50 = in6[50];
    assign x6_51 = in6[51];
    assign x6_52 = in6[52];
    assign x6_53 = in6[53];
    assign x6_54 = in6[54];
    assign x6_55 = in6[55];
    assign x6_56 = in6[56];
    assign x6_57 = in6[57];
    assign x6_58 = in6[58];
    assign x6_59 = in6[59];
    assign x6_60 = in6[60];
    assign x6_61 = in6[61];
    assign x6_62 = in6[62];
    assign x6_63 = in6[63];
    assign x6_64 = in6[64];
    assign x6_65 = in6[65];
    assign x6_66 = in6[66];
    assign x6_67 = in6[67];
    assign x6_68 = in6[68];
    assign x6_69 = in6[69];
    assign x6_70 = in6[70];
    wire x7_0;
    wire x7_1;
    wire x7_2;
    wire x7_3;
    wire x7_4;
    wire x7_5;
    wire x7_6;
    wire x7_7;
    wire x7_8;
    wire x7_9;
    wire x7_10;
    wire x7_11;
    wire x7_12;
    wire x7_13;
    wire x7_14;
    wire x7_15;
    wire x7_16;
    wire x7_17;
    wire x7_18;
    wire x7_19;
    wire x7_20;
    wire x7_21;
    wire x7_22;
    wire x7_23;
    wire x7_24;
    wire x7_25;
    wire x7_26;
    wire x7_27;
    wire x7_28;
    wire x7_29;
    wire x7_30;
    wire x7_31;
    wire x7_32;
    wire x7_33;
    wire x7_34;
    wire x7_35;
    wire x7_36;
    wire x7_37;
    wire x7_38;
    wire x7_39;
    wire x7_40;
    wire x7_41;
    wire x7_42;
    wire x7_43;
    wire x7_44;
    wire x7_45;
    wire x7_46;
    wire x7_47;
    wire x7_48;
    wire x7_49;
    wire x7_50;
    wire x7_51;
    wire x7_52;
    wire x7_53;
    wire x7_54;
    wire x7_55;
    wire x7_56;
    wire x7_57;
    wire x7_58;
    wire x7_59;
    wire x7_60;
    wire x7_61;
    wire x7_62;
    wire x7_63;
    wire x7_64;
    wire x7_65;
    wire x7_66;
    wire x7_67;
    wire x7_68;
    wire x7_69;
    wire x7_70;
    assign x7_0 = in7[0];
    assign x7_1 = in7[1];
    assign x7_2 = in7[2];
    assign x7_3 = in7[3];
    assign x7_4 = in7[4];
    assign x7_5 = in7[5];
    assign x7_6 = in7[6];
    assign x7_7 = in7[7];
    assign x7_8 = in7[8];
    assign x7_9 = in7[9];
    assign x7_10 = in7[10];
    assign x7_11 = in7[11];
    assign x7_12 = in7[12];
    assign x7_13 = in7[13];
    assign x7_14 = in7[14];
    assign x7_15 = in7[15];
    assign x7_16 = in7[16];
    assign x7_17 = in7[17];
    assign x7_18 = in7[18];
    assign x7_19 = in7[19];
    assign x7_20 = in7[20];
    assign x7_21 = in7[21];
    assign x7_22 = in7[22];
    assign x7_23 = in7[23];
    assign x7_24 = in7[24];
    assign x7_25 = in7[25];
    assign x7_26 = in7[26];
    assign x7_27 = in7[27];
    assign x7_28 = in7[28];
    assign x7_29 = in7[29];
    assign x7_30 = in7[30];
    assign x7_31 = in7[31];
    assign x7_32 = in7[32];
    assign x7_33 = in7[33];
    assign x7_34 = in7[34];
    assign x7_35 = in7[35];
    assign x7_36 = in7[36];
    assign x7_37 = in7[37];
    assign x7_38 = in7[38];
    assign x7_39 = in7[39];
    assign x7_40 = in7[40];
    assign x7_41 = in7[41];
    assign x7_42 = in7[42];
    assign x7_43 = in7[43];
    assign x7_44 = in7[44];
    assign x7_45 = in7[45];
    assign x7_46 = in7[46];
    assign x7_47 = in7[47];
    assign x7_48 = in7[48];
    assign x7_49 = in7[49];
    assign x7_50 = in7[50];
    assign x7_51 = in7[51];
    assign x7_52 = in7[52];
    assign x7_53 = in7[53];
    assign x7_54 = in7[54];
    assign x7_55 = in7[55];
    assign x7_56 = in7[56];
    assign x7_57 = in7[57];
    assign x7_58 = in7[58];
    assign x7_59 = in7[59];
    assign x7_60 = in7[60];
    assign x7_61 = in7[61];
    assign x7_62 = in7[62];
    assign x7_63 = in7[63];
    assign x7_64 = in7[64];
    assign x7_65 = in7[65];
    assign x7_66 = in7[66];
    assign x7_67 = in7[67];
    assign x7_68 = in7[68];
    assign x7_69 = in7[69];
    assign x7_70 = in7[70];
    wire x8_0;
    wire x8_1;
    wire x8_2;
    wire x8_3;
    wire x8_4;
    wire x8_5;
    wire x8_6;
    wire x8_7;
    wire x8_8;
    wire x8_9;
    wire x8_10;
    wire x8_11;
    wire x8_12;
    wire x8_13;
    wire x8_14;
    wire x8_15;
    wire x8_16;
    wire x8_17;
    wire x8_18;
    wire x8_19;
    wire x8_20;
    wire x8_21;
    wire x8_22;
    wire x8_23;
    wire x8_24;
    wire x8_25;
    wire x8_26;
    wire x8_27;
    wire x8_28;
    wire x8_29;
    wire x8_30;
    wire x8_31;
    wire x8_32;
    wire x8_33;
    wire x8_34;
    wire x8_35;
    wire x8_36;
    wire x8_37;
    wire x8_38;
    wire x8_39;
    wire x8_40;
    wire x8_41;
    wire x8_42;
    wire x8_43;
    wire x8_44;
    wire x8_45;
    wire x8_46;
    wire x8_47;
    wire x8_48;
    wire x8_49;
    wire x8_50;
    wire x8_51;
    wire x8_52;
    wire x8_53;
    wire x8_54;
    wire x8_55;
    wire x8_56;
    wire x8_57;
    wire x8_58;
    wire x8_59;
    wire x8_60;
    wire x8_61;
    wire x8_62;
    wire x8_63;
    wire x8_64;
    wire x8_65;
    wire x8_66;
    wire x8_67;
    wire x8_68;
    wire x8_69;
    wire x8_70;
    assign x8_0 = in8[0];
    assign x8_1 = in8[1];
    assign x8_2 = in8[2];
    assign x8_3 = in8[3];
    assign x8_4 = in8[4];
    assign x8_5 = in8[5];
    assign x8_6 = in8[6];
    assign x8_7 = in8[7];
    assign x8_8 = in8[8];
    assign x8_9 = in8[9];
    assign x8_10 = in8[10];
    assign x8_11 = in8[11];
    assign x8_12 = in8[12];
    assign x8_13 = in8[13];
    assign x8_14 = in8[14];
    assign x8_15 = in8[15];
    assign x8_16 = in8[16];
    assign x8_17 = in8[17];
    assign x8_18 = in8[18];
    assign x8_19 = in8[19];
    assign x8_20 = in8[20];
    assign x8_21 = in8[21];
    assign x8_22 = in8[22];
    assign x8_23 = in8[23];
    assign x8_24 = in8[24];
    assign x8_25 = in8[25];
    assign x8_26 = in8[26];
    assign x8_27 = in8[27];
    assign x8_28 = in8[28];
    assign x8_29 = in8[29];
    assign x8_30 = in8[30];
    assign x8_31 = in8[31];
    assign x8_32 = in8[32];
    assign x8_33 = in8[33];
    assign x8_34 = in8[34];
    assign x8_35 = in8[35];
    assign x8_36 = in8[36];
    assign x8_37 = in8[37];
    assign x8_38 = in8[38];
    assign x8_39 = in8[39];
    assign x8_40 = in8[40];
    assign x8_41 = in8[41];
    assign x8_42 = in8[42];
    assign x8_43 = in8[43];
    assign x8_44 = in8[44];
    assign x8_45 = in8[45];
    assign x8_46 = in8[46];
    assign x8_47 = in8[47];
    assign x8_48 = in8[48];
    assign x8_49 = in8[49];
    assign x8_50 = in8[50];
    assign x8_51 = in8[51];
    assign x8_52 = in8[52];
    assign x8_53 = in8[53];
    assign x8_54 = in8[54];
    assign x8_55 = in8[55];
    assign x8_56 = in8[56];
    assign x8_57 = in8[57];
    assign x8_58 = in8[58];
    assign x8_59 = in8[59];
    assign x8_60 = in8[60];
    assign x8_61 = in8[61];
    assign x8_62 = in8[62];
    assign x8_63 = in8[63];
    assign x8_64 = in8[64];
    assign x8_65 = in8[65];
    assign x8_66 = in8[66];
    assign x8_67 = in8[67];
    assign x8_68 = in8[68];
    assign x8_69 = in8[69];
    assign x8_70 = in8[70];
    wire x9_0;
    wire x9_1;
    wire x9_2;
    wire x9_3;
    wire x9_4;
    wire x9_5;
    wire x9_6;
    wire x9_7;
    wire x9_8;
    wire x9_9;
    wire x9_10;
    wire x9_11;
    wire x9_12;
    wire x9_13;
    wire x9_14;
    wire x9_15;
    wire x9_16;
    wire x9_17;
    wire x9_18;
    wire x9_19;
    wire x9_20;
    wire x9_21;
    wire x9_22;
    wire x9_23;
    wire x9_24;
    wire x9_25;
    wire x9_26;
    wire x9_27;
    wire x9_28;
    wire x9_29;
    wire x9_30;
    wire x9_31;
    wire x9_32;
    wire x9_33;
    wire x9_34;
    wire x9_35;
    wire x9_36;
    wire x9_37;
    wire x9_38;
    wire x9_39;
    wire x9_40;
    wire x9_41;
    wire x9_42;
    wire x9_43;
    wire x9_44;
    wire x9_45;
    wire x9_46;
    wire x9_47;
    wire x9_48;
    wire x9_49;
    wire x9_50;
    wire x9_51;
    wire x9_52;
    wire x9_53;
    wire x9_54;
    wire x9_55;
    wire x9_56;
    wire x9_57;
    wire x9_58;
    wire x9_59;
    wire x9_60;
    wire x9_61;
    wire x9_62;
    wire x9_63;
    wire x9_64;
    wire x9_65;
    wire x9_66;
    wire x9_67;
    wire x9_68;
    wire x9_69;
    wire x9_70;
    assign x9_0 = in9[0];
    assign x9_1 = in9[1];
    assign x9_2 = in9[2];
    assign x9_3 = in9[3];
    assign x9_4 = in9[4];
    assign x9_5 = in9[5];
    assign x9_6 = in9[6];
    assign x9_7 = in9[7];
    assign x9_8 = in9[8];
    assign x9_9 = in9[9];
    assign x9_10 = in9[10];
    assign x9_11 = in9[11];
    assign x9_12 = in9[12];
    assign x9_13 = in9[13];
    assign x9_14 = in9[14];
    assign x9_15 = in9[15];
    assign x9_16 = in9[16];
    assign x9_17 = in9[17];
    assign x9_18 = in9[18];
    assign x9_19 = in9[19];
    assign x9_20 = in9[20];
    assign x9_21 = in9[21];
    assign x9_22 = in9[22];
    assign x9_23 = in9[23];
    assign x9_24 = in9[24];
    assign x9_25 = in9[25];
    assign x9_26 = in9[26];
    assign x9_27 = in9[27];
    assign x9_28 = in9[28];
    assign x9_29 = in9[29];
    assign x9_30 = in9[30];
    assign x9_31 = in9[31];
    assign x9_32 = in9[32];
    assign x9_33 = in9[33];
    assign x9_34 = in9[34];
    assign x9_35 = in9[35];
    assign x9_36 = in9[36];
    assign x9_37 = in9[37];
    assign x9_38 = in9[38];
    assign x9_39 = in9[39];
    assign x9_40 = in9[40];
    assign x9_41 = in9[41];
    assign x9_42 = in9[42];
    assign x9_43 = in9[43];
    assign x9_44 = in9[44];
    assign x9_45 = in9[45];
    assign x9_46 = in9[46];
    assign x9_47 = in9[47];
    assign x9_48 = in9[48];
    assign x9_49 = in9[49];
    assign x9_50 = in9[50];
    assign x9_51 = in9[51];
    assign x9_52 = in9[52];
    assign x9_53 = in9[53];
    assign x9_54 = in9[54];
    assign x9_55 = in9[55];
    assign x9_56 = in9[56];
    assign x9_57 = in9[57];
    assign x9_58 = in9[58];
    assign x9_59 = in9[59];
    assign x9_60 = in9[60];
    assign x9_61 = in9[61];
    assign x9_62 = in9[62];
    assign x9_63 = in9[63];
    assign x9_64 = in9[64];
    assign x9_65 = in9[65];
    assign x9_66 = in9[66];
    assign x9_67 = in9[67];
    assign x9_68 = in9[68];
    assign x9_69 = in9[69];
    assign x9_70 = in9[70];
    wire x10_0;
    wire x10_1;
    wire x10_2;
    wire x10_3;
    wire x10_4;
    wire x10_5;
    wire x10_6;
    wire x10_7;
    wire x10_8;
    wire x10_9;
    wire x10_10;
    wire x10_11;
    wire x10_12;
    wire x10_13;
    wire x10_14;
    wire x10_15;
    wire x10_16;
    wire x10_17;
    wire x10_18;
    wire x10_19;
    wire x10_20;
    wire x10_21;
    wire x10_22;
    wire x10_23;
    wire x10_24;
    wire x10_25;
    wire x10_26;
    wire x10_27;
    wire x10_28;
    wire x10_29;
    wire x10_30;
    wire x10_31;
    wire x10_32;
    wire x10_33;
    wire x10_34;
    wire x10_35;
    wire x10_36;
    wire x10_37;
    wire x10_38;
    wire x10_39;
    wire x10_40;
    wire x10_41;
    wire x10_42;
    wire x10_43;
    wire x10_44;
    wire x10_45;
    wire x10_46;
    wire x10_47;
    wire x10_48;
    wire x10_49;
    wire x10_50;
    wire x10_51;
    wire x10_52;
    wire x10_53;
    wire x10_54;
    wire x10_55;
    wire x10_56;
    wire x10_57;
    wire x10_58;
    wire x10_59;
    wire x10_60;
    wire x10_61;
    wire x10_62;
    wire x10_63;
    wire x10_64;
    wire x10_65;
    wire x10_66;
    wire x10_67;
    wire x10_68;
    wire x10_69;
    wire x10_70;
    assign x10_0 = in10[0];
    assign x10_1 = in10[1];
    assign x10_2 = in10[2];
    assign x10_3 = in10[3];
    assign x10_4 = in10[4];
    assign x10_5 = in10[5];
    assign x10_6 = in10[6];
    assign x10_7 = in10[7];
    assign x10_8 = in10[8];
    assign x10_9 = in10[9];
    assign x10_10 = in10[10];
    assign x10_11 = in10[11];
    assign x10_12 = in10[12];
    assign x10_13 = in10[13];
    assign x10_14 = in10[14];
    assign x10_15 = in10[15];
    assign x10_16 = in10[16];
    assign x10_17 = in10[17];
    assign x10_18 = in10[18];
    assign x10_19 = in10[19];
    assign x10_20 = in10[20];
    assign x10_21 = in10[21];
    assign x10_22 = in10[22];
    assign x10_23 = in10[23];
    assign x10_24 = in10[24];
    assign x10_25 = in10[25];
    assign x10_26 = in10[26];
    assign x10_27 = in10[27];
    assign x10_28 = in10[28];
    assign x10_29 = in10[29];
    assign x10_30 = in10[30];
    assign x10_31 = in10[31];
    assign x10_32 = in10[32];
    assign x10_33 = in10[33];
    assign x10_34 = in10[34];
    assign x10_35 = in10[35];
    assign x10_36 = in10[36];
    assign x10_37 = in10[37];
    assign x10_38 = in10[38];
    assign x10_39 = in10[39];
    assign x10_40 = in10[40];
    assign x10_41 = in10[41];
    assign x10_42 = in10[42];
    assign x10_43 = in10[43];
    assign x10_44 = in10[44];
    assign x10_45 = in10[45];
    assign x10_46 = in10[46];
    assign x10_47 = in10[47];
    assign x10_48 = in10[48];
    assign x10_49 = in10[49];
    assign x10_50 = in10[50];
    assign x10_51 = in10[51];
    assign x10_52 = in10[52];
    assign x10_53 = in10[53];
    assign x10_54 = in10[54];
    assign x10_55 = in10[55];
    assign x10_56 = in10[56];
    assign x10_57 = in10[57];
    assign x10_58 = in10[58];
    assign x10_59 = in10[59];
    assign x10_60 = in10[60];
    assign x10_61 = in10[61];
    assign x10_62 = in10[62];
    assign x10_63 = in10[63];
    assign x10_64 = in10[64];
    assign x10_65 = in10[65];
    assign x10_66 = in10[66];
    assign x10_67 = in10[67];
    assign x10_68 = in10[68];
    assign x10_69 = in10[69];
    assign x10_70 = in10[70];
    wire x11_0;
    wire x11_1;
    wire x11_2;
    wire x11_3;
    wire x11_4;
    wire x11_5;
    wire x11_6;
    wire x11_7;
    wire x11_8;
    wire x11_9;
    wire x11_10;
    wire x11_11;
    wire x11_12;
    wire x11_13;
    wire x11_14;
    wire x11_15;
    wire x11_16;
    wire x11_17;
    wire x11_18;
    wire x11_19;
    wire x11_20;
    wire x11_21;
    wire x11_22;
    wire x11_23;
    wire x11_24;
    wire x11_25;
    wire x11_26;
    wire x11_27;
    wire x11_28;
    wire x11_29;
    wire x11_30;
    wire x11_31;
    wire x11_32;
    wire x11_33;
    wire x11_34;
    wire x11_35;
    wire x11_36;
    wire x11_37;
    wire x11_38;
    wire x11_39;
    wire x11_40;
    wire x11_41;
    wire x11_42;
    wire x11_43;
    wire x11_44;
    wire x11_45;
    wire x11_46;
    wire x11_47;
    wire x11_48;
    wire x11_49;
    wire x11_50;
    wire x11_51;
    wire x11_52;
    wire x11_53;
    wire x11_54;
    wire x11_55;
    wire x11_56;
    wire x11_57;
    wire x11_58;
    wire x11_59;
    wire x11_60;
    wire x11_61;
    wire x11_62;
    wire x11_63;
    wire x11_64;
    wire x11_65;
    wire x11_66;
    wire x11_67;
    wire x11_68;
    wire x11_69;
    wire x11_70;
    assign x11_0 = in11[0];
    assign x11_1 = in11[1];
    assign x11_2 = in11[2];
    assign x11_3 = in11[3];
    assign x11_4 = in11[4];
    assign x11_5 = in11[5];
    assign x11_6 = in11[6];
    assign x11_7 = in11[7];
    assign x11_8 = in11[8];
    assign x11_9 = in11[9];
    assign x11_10 = in11[10];
    assign x11_11 = in11[11];
    assign x11_12 = in11[12];
    assign x11_13 = in11[13];
    assign x11_14 = in11[14];
    assign x11_15 = in11[15];
    assign x11_16 = in11[16];
    assign x11_17 = in11[17];
    assign x11_18 = in11[18];
    assign x11_19 = in11[19];
    assign x11_20 = in11[20];
    assign x11_21 = in11[21];
    assign x11_22 = in11[22];
    assign x11_23 = in11[23];
    assign x11_24 = in11[24];
    assign x11_25 = in11[25];
    assign x11_26 = in11[26];
    assign x11_27 = in11[27];
    assign x11_28 = in11[28];
    assign x11_29 = in11[29];
    assign x11_30 = in11[30];
    assign x11_31 = in11[31];
    assign x11_32 = in11[32];
    assign x11_33 = in11[33];
    assign x11_34 = in11[34];
    assign x11_35 = in11[35];
    assign x11_36 = in11[36];
    assign x11_37 = in11[37];
    assign x11_38 = in11[38];
    assign x11_39 = in11[39];
    assign x11_40 = in11[40];
    assign x11_41 = in11[41];
    assign x11_42 = in11[42];
    assign x11_43 = in11[43];
    assign x11_44 = in11[44];
    assign x11_45 = in11[45];
    assign x11_46 = in11[46];
    assign x11_47 = in11[47];
    assign x11_48 = in11[48];
    assign x11_49 = in11[49];
    assign x11_50 = in11[50];
    assign x11_51 = in11[51];
    assign x11_52 = in11[52];
    assign x11_53 = in11[53];
    assign x11_54 = in11[54];
    assign x11_55 = in11[55];
    assign x11_56 = in11[56];
    assign x11_57 = in11[57];
    assign x11_58 = in11[58];
    assign x11_59 = in11[59];
    assign x11_60 = in11[60];
    assign x11_61 = in11[61];
    assign x11_62 = in11[62];
    assign x11_63 = in11[63];
    assign x11_64 = in11[64];
    assign x11_65 = in11[65];
    assign x11_66 = in11[66];
    assign x11_67 = in11[67];
    assign x11_68 = in11[68];
    assign x11_69 = in11[69];
    assign x11_70 = in11[70];
    wire x12_0;
    wire x12_1;
    wire x12_2;
    wire x12_3;
    wire x12_4;
    wire x12_5;
    wire x12_6;
    wire x12_7;
    wire x12_8;
    wire x12_9;
    wire x12_10;
    wire x12_11;
    wire x12_12;
    wire x12_13;
    wire x12_14;
    wire x12_15;
    wire x12_16;
    wire x12_17;
    wire x12_18;
    wire x12_19;
    wire x12_20;
    wire x12_21;
    wire x12_22;
    wire x12_23;
    wire x12_24;
    wire x12_25;
    wire x12_26;
    wire x12_27;
    wire x12_28;
    wire x12_29;
    wire x12_30;
    wire x12_31;
    wire x12_32;
    wire x12_33;
    wire x12_34;
    wire x12_35;
    wire x12_36;
    wire x12_37;
    wire x12_38;
    wire x12_39;
    wire x12_40;
    wire x12_41;
    wire x12_42;
    wire x12_43;
    wire x12_44;
    wire x12_45;
    wire x12_46;
    wire x12_47;
    wire x12_48;
    wire x12_49;
    wire x12_50;
    wire x12_51;
    wire x12_52;
    wire x12_53;
    wire x12_54;
    wire x12_55;
    wire x12_56;
    wire x12_57;
    wire x12_58;
    wire x12_59;
    wire x12_60;
    wire x12_61;
    wire x12_62;
    wire x12_63;
    wire x12_64;
    wire x12_65;
    wire x12_66;
    wire x12_67;
    wire x12_68;
    wire x12_69;
    wire x12_70;
    assign x12_0 = in12[0];
    assign x12_1 = in12[1];
    assign x12_2 = in12[2];
    assign x12_3 = in12[3];
    assign x12_4 = in12[4];
    assign x12_5 = in12[5];
    assign x12_6 = in12[6];
    assign x12_7 = in12[7];
    assign x12_8 = in12[8];
    assign x12_9 = in12[9];
    assign x12_10 = in12[10];
    assign x12_11 = in12[11];
    assign x12_12 = in12[12];
    assign x12_13 = in12[13];
    assign x12_14 = in12[14];
    assign x12_15 = in12[15];
    assign x12_16 = in12[16];
    assign x12_17 = in12[17];
    assign x12_18 = in12[18];
    assign x12_19 = in12[19];
    assign x12_20 = in12[20];
    assign x12_21 = in12[21];
    assign x12_22 = in12[22];
    assign x12_23 = in12[23];
    assign x12_24 = in12[24];
    assign x12_25 = in12[25];
    assign x12_26 = in12[26];
    assign x12_27 = in12[27];
    assign x12_28 = in12[28];
    assign x12_29 = in12[29];
    assign x12_30 = in12[30];
    assign x12_31 = in12[31];
    assign x12_32 = in12[32];
    assign x12_33 = in12[33];
    assign x12_34 = in12[34];
    assign x12_35 = in12[35];
    assign x12_36 = in12[36];
    assign x12_37 = in12[37];
    assign x12_38 = in12[38];
    assign x12_39 = in12[39];
    assign x12_40 = in12[40];
    assign x12_41 = in12[41];
    assign x12_42 = in12[42];
    assign x12_43 = in12[43];
    assign x12_44 = in12[44];
    assign x12_45 = in12[45];
    assign x12_46 = in12[46];
    assign x12_47 = in12[47];
    assign x12_48 = in12[48];
    assign x12_49 = in12[49];
    assign x12_50 = in12[50];
    assign x12_51 = in12[51];
    assign x12_52 = in12[52];
    assign x12_53 = in12[53];
    assign x12_54 = in12[54];
    assign x12_55 = in12[55];
    assign x12_56 = in12[56];
    assign x12_57 = in12[57];
    assign x12_58 = in12[58];
    assign x12_59 = in12[59];
    assign x12_60 = in12[60];
    assign x12_61 = in12[61];
    assign x12_62 = in12[62];
    assign x12_63 = in12[63];
    assign x12_64 = in12[64];
    assign x12_65 = in12[65];
    assign x12_66 = in12[66];
    assign x12_67 = in12[67];
    assign x12_68 = in12[68];
    assign x12_69 = in12[69];
    assign x12_70 = in12[70];
    wire x13_0;
    wire x13_1;
    wire x13_2;
    wire x13_3;
    wire x13_4;
    wire x13_5;
    wire x13_6;
    wire x13_7;
    wire x13_8;
    wire x13_9;
    wire x13_10;
    wire x13_11;
    wire x13_12;
    wire x13_13;
    wire x13_14;
    wire x13_15;
    wire x13_16;
    wire x13_17;
    wire x13_18;
    wire x13_19;
    wire x13_20;
    wire x13_21;
    wire x13_22;
    wire x13_23;
    wire x13_24;
    wire x13_25;
    wire x13_26;
    wire x13_27;
    wire x13_28;
    wire x13_29;
    wire x13_30;
    wire x13_31;
    wire x13_32;
    wire x13_33;
    wire x13_34;
    wire x13_35;
    wire x13_36;
    wire x13_37;
    wire x13_38;
    wire x13_39;
    wire x13_40;
    wire x13_41;
    wire x13_42;
    wire x13_43;
    wire x13_44;
    wire x13_45;
    wire x13_46;
    wire x13_47;
    wire x13_48;
    wire x13_49;
    wire x13_50;
    wire x13_51;
    wire x13_52;
    wire x13_53;
    wire x13_54;
    wire x13_55;
    wire x13_56;
    wire x13_57;
    wire x13_58;
    wire x13_59;
    wire x13_60;
    wire x13_61;
    wire x13_62;
    wire x13_63;
    wire x13_64;
    wire x13_65;
    wire x13_66;
    wire x13_67;
    wire x13_68;
    wire x13_69;
    wire x13_70;
    assign x13_0 = in13[0];
    assign x13_1 = in13[1];
    assign x13_2 = in13[2];
    assign x13_3 = in13[3];
    assign x13_4 = in13[4];
    assign x13_5 = in13[5];
    assign x13_6 = in13[6];
    assign x13_7 = in13[7];
    assign x13_8 = in13[8];
    assign x13_9 = in13[9];
    assign x13_10 = in13[10];
    assign x13_11 = in13[11];
    assign x13_12 = in13[12];
    assign x13_13 = in13[13];
    assign x13_14 = in13[14];
    assign x13_15 = in13[15];
    assign x13_16 = in13[16];
    assign x13_17 = in13[17];
    assign x13_18 = in13[18];
    assign x13_19 = in13[19];
    assign x13_20 = in13[20];
    assign x13_21 = in13[21];
    assign x13_22 = in13[22];
    assign x13_23 = in13[23];
    assign x13_24 = in13[24];
    assign x13_25 = in13[25];
    assign x13_26 = in13[26];
    assign x13_27 = in13[27];
    assign x13_28 = in13[28];
    assign x13_29 = in13[29];
    assign x13_30 = in13[30];
    assign x13_31 = in13[31];
    assign x13_32 = in13[32];
    assign x13_33 = in13[33];
    assign x13_34 = in13[34];
    assign x13_35 = in13[35];
    assign x13_36 = in13[36];
    assign x13_37 = in13[37];
    assign x13_38 = in13[38];
    assign x13_39 = in13[39];
    assign x13_40 = in13[40];
    assign x13_41 = in13[41];
    assign x13_42 = in13[42];
    assign x13_43 = in13[43];
    assign x13_44 = in13[44];
    assign x13_45 = in13[45];
    assign x13_46 = in13[46];
    assign x13_47 = in13[47];
    assign x13_48 = in13[48];
    assign x13_49 = in13[49];
    assign x13_50 = in13[50];
    assign x13_51 = in13[51];
    assign x13_52 = in13[52];
    assign x13_53 = in13[53];
    assign x13_54 = in13[54];
    assign x13_55 = in13[55];
    assign x13_56 = in13[56];
    assign x13_57 = in13[57];
    assign x13_58 = in13[58];
    assign x13_59 = in13[59];
    assign x13_60 = in13[60];
    assign x13_61 = in13[61];
    assign x13_62 = in13[62];
    assign x13_63 = in13[63];
    assign x13_64 = in13[64];
    assign x13_65 = in13[65];
    assign x13_66 = in13[66];
    assign x13_67 = in13[67];
    assign x13_68 = in13[68];
    assign x13_69 = in13[69];
    assign x13_70 = in13[70];
    wire x14_0;
    wire x14_1;
    wire x14_2;
    wire x14_3;
    wire x14_4;
    wire x14_5;
    wire x14_6;
    wire x14_7;
    wire x14_8;
    wire x14_9;
    wire x14_10;
    wire x14_11;
    wire x14_12;
    wire x14_13;
    wire x14_14;
    wire x14_15;
    wire x14_16;
    wire x14_17;
    wire x14_18;
    wire x14_19;
    wire x14_20;
    wire x14_21;
    wire x14_22;
    wire x14_23;
    wire x14_24;
    wire x14_25;
    wire x14_26;
    wire x14_27;
    wire x14_28;
    wire x14_29;
    wire x14_30;
    wire x14_31;
    wire x14_32;
    wire x14_33;
    wire x14_34;
    wire x14_35;
    wire x14_36;
    wire x14_37;
    wire x14_38;
    wire x14_39;
    wire x14_40;
    wire x14_41;
    wire x14_42;
    wire x14_43;
    wire x14_44;
    wire x14_45;
    wire x14_46;
    wire x14_47;
    wire x14_48;
    wire x14_49;
    wire x14_50;
    wire x14_51;
    wire x14_52;
    wire x14_53;
    wire x14_54;
    wire x14_55;
    wire x14_56;
    wire x14_57;
    wire x14_58;
    wire x14_59;
    wire x14_60;
    wire x14_61;
    wire x14_62;
    wire x14_63;
    wire x14_64;
    wire x14_65;
    wire x14_66;
    wire x14_67;
    wire x14_68;
    wire x14_69;
    wire x14_70;
    assign x14_0 = in14[0];
    assign x14_1 = in14[1];
    assign x14_2 = in14[2];
    assign x14_3 = in14[3];
    assign x14_4 = in14[4];
    assign x14_5 = in14[5];
    assign x14_6 = in14[6];
    assign x14_7 = in14[7];
    assign x14_8 = in14[8];
    assign x14_9 = in14[9];
    assign x14_10 = in14[10];
    assign x14_11 = in14[11];
    assign x14_12 = in14[12];
    assign x14_13 = in14[13];
    assign x14_14 = in14[14];
    assign x14_15 = in14[15];
    assign x14_16 = in14[16];
    assign x14_17 = in14[17];
    assign x14_18 = in14[18];
    assign x14_19 = in14[19];
    assign x14_20 = in14[20];
    assign x14_21 = in14[21];
    assign x14_22 = in14[22];
    assign x14_23 = in14[23];
    assign x14_24 = in14[24];
    assign x14_25 = in14[25];
    assign x14_26 = in14[26];
    assign x14_27 = in14[27];
    assign x14_28 = in14[28];
    assign x14_29 = in14[29];
    assign x14_30 = in14[30];
    assign x14_31 = in14[31];
    assign x14_32 = in14[32];
    assign x14_33 = in14[33];
    assign x14_34 = in14[34];
    assign x14_35 = in14[35];
    assign x14_36 = in14[36];
    assign x14_37 = in14[37];
    assign x14_38 = in14[38];
    assign x14_39 = in14[39];
    assign x14_40 = in14[40];
    assign x14_41 = in14[41];
    assign x14_42 = in14[42];
    assign x14_43 = in14[43];
    assign x14_44 = in14[44];
    assign x14_45 = in14[45];
    assign x14_46 = in14[46];
    assign x14_47 = in14[47];
    assign x14_48 = in14[48];
    assign x14_49 = in14[49];
    assign x14_50 = in14[50];
    assign x14_51 = in14[51];
    assign x14_52 = in14[52];
    assign x14_53 = in14[53];
    assign x14_54 = in14[54];
    assign x14_55 = in14[55];
    assign x14_56 = in14[56];
    assign x14_57 = in14[57];
    assign x14_58 = in14[58];
    assign x14_59 = in14[59];
    assign x14_60 = in14[60];
    assign x14_61 = in14[61];
    assign x14_62 = in14[62];
    assign x14_63 = in14[63];
    assign x14_64 = in14[64];
    assign x14_65 = in14[65];
    assign x14_66 = in14[66];
    assign x14_67 = in14[67];
    assign x14_68 = in14[68];
    assign x14_69 = in14[69];
    assign x14_70 = in14[70];
    wire x15_0;
    wire x15_1;
    wire x15_2;
    wire x15_3;
    wire x15_4;
    wire x15_5;
    wire x15_6;
    wire x15_7;
    wire x15_8;
    wire x15_9;
    wire x15_10;
    wire x15_11;
    wire x15_12;
    wire x15_13;
    wire x15_14;
    wire x15_15;
    wire x15_16;
    wire x15_17;
    wire x15_18;
    wire x15_19;
    wire x15_20;
    wire x15_21;
    wire x15_22;
    wire x15_23;
    wire x15_24;
    wire x15_25;
    wire x15_26;
    wire x15_27;
    wire x15_28;
    wire x15_29;
    wire x15_30;
    wire x15_31;
    wire x15_32;
    wire x15_33;
    wire x15_34;
    wire x15_35;
    wire x15_36;
    wire x15_37;
    wire x15_38;
    wire x15_39;
    wire x15_40;
    wire x15_41;
    wire x15_42;
    wire x15_43;
    wire x15_44;
    wire x15_45;
    wire x15_46;
    wire x15_47;
    wire x15_48;
    wire x15_49;
    wire x15_50;
    wire x15_51;
    wire x15_52;
    wire x15_53;
    wire x15_54;
    wire x15_55;
    wire x15_56;
    wire x15_57;
    wire x15_58;
    wire x15_59;
    wire x15_60;
    wire x15_61;
    wire x15_62;
    wire x15_63;
    wire x15_64;
    wire x15_65;
    wire x15_66;
    wire x15_67;
    wire x15_68;
    wire x15_69;
    wire x15_70;
    assign x15_0 = in15[0];
    assign x15_1 = in15[1];
    assign x15_2 = in15[2];
    assign x15_3 = in15[3];
    assign x15_4 = in15[4];
    assign x15_5 = in15[5];
    assign x15_6 = in15[6];
    assign x15_7 = in15[7];
    assign x15_8 = in15[8];
    assign x15_9 = in15[9];
    assign x15_10 = in15[10];
    assign x15_11 = in15[11];
    assign x15_12 = in15[12];
    assign x15_13 = in15[13];
    assign x15_14 = in15[14];
    assign x15_15 = in15[15];
    assign x15_16 = in15[16];
    assign x15_17 = in15[17];
    assign x15_18 = in15[18];
    assign x15_19 = in15[19];
    assign x15_20 = in15[20];
    assign x15_21 = in15[21];
    assign x15_22 = in15[22];
    assign x15_23 = in15[23];
    assign x15_24 = in15[24];
    assign x15_25 = in15[25];
    assign x15_26 = in15[26];
    assign x15_27 = in15[27];
    assign x15_28 = in15[28];
    assign x15_29 = in15[29];
    assign x15_30 = in15[30];
    assign x15_31 = in15[31];
    assign x15_32 = in15[32];
    assign x15_33 = in15[33];
    assign x15_34 = in15[34];
    assign x15_35 = in15[35];
    assign x15_36 = in15[36];
    assign x15_37 = in15[37];
    assign x15_38 = in15[38];
    assign x15_39 = in15[39];
    assign x15_40 = in15[40];
    assign x15_41 = in15[41];
    assign x15_42 = in15[42];
    assign x15_43 = in15[43];
    assign x15_44 = in15[44];
    assign x15_45 = in15[45];
    assign x15_46 = in15[46];
    assign x15_47 = in15[47];
    assign x15_48 = in15[48];
    assign x15_49 = in15[49];
    assign x15_50 = in15[50];
    assign x15_51 = in15[51];
    assign x15_52 = in15[52];
    assign x15_53 = in15[53];
    assign x15_54 = in15[54];
    assign x15_55 = in15[55];
    assign x15_56 = in15[56];
    assign x15_57 = in15[57];
    assign x15_58 = in15[58];
    assign x15_59 = in15[59];
    assign x15_60 = in15[60];
    assign x15_61 = in15[61];
    assign x15_62 = in15[62];
    assign x15_63 = in15[63];
    assign x15_64 = in15[64];
    assign x15_65 = in15[65];
    assign x15_66 = in15[66];
    assign x15_67 = in15[67];
    assign x15_68 = in15[68];
    assign x15_69 = in15[69];
    assign x15_70 = in15[70];
    wire w287;
    wire w288;
    wire w289;
    wire w290;
    wire w291;
    wire w292;
    wire w293;
    wire w294;
    wire w295;
    wire w296;
    wire w297;
    wire w298;
    wire w299;
    wire w300;
    wire w301;
    wire w302;
    wire w303;
    wire w304;
    wire w305;
    wire w306;
    wire w307;
    wire w308;
    wire w309;
    wire w310;
    wire w311;
    wire w312;
    wire w313;
    wire w314;
    wire w315;
    wire w316;
    wire w317;
    wire w318;
    wire w319;
    wire w320;
    wire w321;
    wire w322;
    wire w323;
    wire w324;
    wire w325;
    wire w326;
    wire w327;
    wire w328;
    wire w329;
    wire w330;
    wire w331;
    wire w332;
    wire w333;
    wire w334;
    wire w335;
    wire w336;
    wire w337;
    wire w338;
    wire w339;
    wire w340;
    wire w341;
    wire w342;
    wire w343;
    wire w344;
    wire w345;
    wire w346;
    wire w347;
    wire w348;
    wire w349;
    wire w350;
    wire w351;
    wire w352;
    wire w353;
    wire w354;
    wire w355;
    wire w356;
    assign out0[0] = w287;
    assign out0[1] = w288;
    assign out0[2] = w289;
    assign out0[3] = w290;
    assign out0[4] = w291;
    assign out0[5] = w292;
    assign out0[6] = w293;
    assign out0[7] = w294;
    assign out0[8] = w295;
    assign out0[9] = w296;
    assign out0[10] = w297;
    assign out0[11] = w298;
    assign out0[12] = w299;
    assign out0[13] = w300;
    assign out0[14] = w301;
    assign out0[15] = w302;
    assign out0[16] = w303;
    assign out0[17] = w304;
    assign out0[18] = w305;
    assign out0[19] = w306;
    assign out0[20] = w307;
    assign out0[21] = w308;
    assign out0[22] = w309;
    assign out0[23] = w310;
    assign out0[24] = w311;
    assign out0[25] = w312;
    assign out0[26] = w313;
    assign out0[27] = w314;
    assign out0[28] = w315;
    assign out0[29] = w316;
    assign out0[30] = w317;
    assign out0[31] = w318;
    assign out0[32] = w319;
    assign out0[33] = w320;
    assign out0[34] = w321;
    assign out0[35] = w322;
    assign out0[36] = w323;
    assign out0[37] = w324;
    assign out0[38] = w325;
    assign out0[39] = w326;
    assign out0[40] = w327;
    assign out0[41] = w328;
    assign out0[42] = w329;
    assign out0[43] = w330;
    assign out0[44] = w331;
    assign out0[45] = w332;
    assign out0[46] = w333;
    assign out0[47] = w334;
    assign out0[48] = w335;
    assign out0[49] = w336;
    assign out0[50] = w337;
    assign out0[51] = w338;
    assign out0[52] = w339;
    assign out0[53] = w340;
    assign out0[54] = w341;
    assign out0[55] = w342;
    assign out0[56] = w343;
    assign out0[57] = w344;
    assign out0[58] = w345;
    assign out0[59] = w346;
    assign out0[60] = w347;
    assign out0[61] = w348;
    assign out0[62] = w349;
    assign out0[63] = w350;
    assign out0[64] = w351;
    assign out0[65] = w352;
    assign out0[66] = w353;
    assign out0[67] = w354;
    assign out0[68] = w355;
    assign out0[69] = w356;
    wire w427;
    wire w428;
    wire w429;
    wire w430;
    wire w431;
    wire w432;
    wire w433;
    wire w434;
    wire w435;
    wire w436;
    wire w437;
    wire w438;
    wire w439;
    wire w440;
    wire w441;
    wire w442;
    wire w443;
    wire w444;
    wire w445;
    wire w446;
    wire w447;
    wire w448;
    wire w449;
    wire w450;
    wire w451;
    wire w452;
    wire w453;
    wire w454;
    wire w455;
    wire w456;
    wire w457;
    wire w458;
    wire w459;
    wire w460;
    wire w461;
    wire w462;
    wire w463;
    wire w464;
    wire w465;
    wire w466;
    wire w467;
    wire w468;
    wire w469;
    wire w470;
    wire w471;
    wire w472;
    wire w473;
    wire w474;
    wire w475;
    wire w476;
    wire w477;
    wire w478;
    wire w479;
    wire w480;
    wire w481;
    wire w482;
    wire w483;
    wire w484;
    wire w485;
    wire w486;
    wire w487;
    wire w488;
    wire w489;
    wire w490;
    wire w491;
    wire w492;
    wire w493;
    wire w494;
    wire w495;
    wire w496;
    assign out1[0] = w427;
    assign out1[1] = w428;
    assign out1[2] = w429;
    assign out1[3] = w430;
    assign out1[4] = w431;
    assign out1[5] = w432;
    assign out1[6] = w433;
    assign out1[7] = w434;
    assign out1[8] = w435;
    assign out1[9] = w436;
    assign out1[10] = w437;
    assign out1[11] = w438;
    assign out1[12] = w439;
    assign out1[13] = w440;
    assign out1[14] = w441;
    assign out1[15] = w442;
    assign out1[16] = w443;
    assign out1[17] = w444;
    assign out1[18] = w445;
    assign out1[19] = w446;
    assign out1[20] = w447;
    assign out1[21] = w448;
    assign out1[22] = w449;
    assign out1[23] = w450;
    assign out1[24] = w451;
    assign out1[25] = w452;
    assign out1[26] = w453;
    assign out1[27] = w454;
    assign out1[28] = w455;
    assign out1[29] = w456;
    assign out1[30] = w457;
    assign out1[31] = w458;
    assign out1[32] = w459;
    assign out1[33] = w460;
    assign out1[34] = w461;
    assign out1[35] = w462;
    assign out1[36] = w463;
    assign out1[37] = w464;
    assign out1[38] = w465;
    assign out1[39] = w466;
    assign out1[40] = w467;
    assign out1[41] = w468;
    assign out1[42] = w469;
    assign out1[43] = w470;
    assign out1[44] = w471;
    assign out1[45] = w472;
    assign out1[46] = w473;
    assign out1[47] = w474;
    assign out1[48] = w475;
    assign out1[49] = w476;
    assign out1[50] = w477;
    assign out1[51] = w478;
    assign out1[52] = w479;
    assign out1[53] = w480;
    assign out1[54] = w481;
    assign out1[55] = w482;
    assign out1[56] = w483;
    assign out1[57] = w484;
    assign out1[58] = w485;
    assign out1[59] = w486;
    assign out1[60] = w487;
    assign out1[61] = w488;
    assign out1[62] = w489;
    assign out1[63] = w490;
    assign out1[64] = w491;
    assign out1[65] = w492;
    assign out1[66] = w493;
    assign out1[67] = w494;
    assign out1[68] = w495;
    assign out1[69] = w496;
    wire w497;
    wire w498;
    wire w499;
    wire w500;
    wire w501;
    wire w502;
    wire w503;
    wire w504;
    wire w505;
    wire w506;
    wire w507;
    wire w508;
    wire w509;
    wire w510;
    wire w511;
    wire w512;
    wire w513;
    wire w514;
    wire w515;
    wire w516;
    wire w517;
    wire w518;
    wire w519;
    wire w520;
    wire w521;
    wire w522;
    wire w523;
    wire w524;
    wire w525;
    wire w526;
    wire w527;
    wire w528;
    wire w529;
    wire w530;
    wire w531;
    wire w532;
    wire w533;
    wire w534;
    wire w535;
    wire w536;
    wire w537;
    wire w538;
    wire w539;
    wire w540;
    wire w541;
    wire w542;
    wire w543;
    wire w544;
    wire w545;
    wire w546;
    wire w547;
    wire w548;
    wire w549;
    wire w550;
    wire w551;
    wire w552;
    wire w553;
    wire w554;
    wire w555;
    wire w556;
    wire w557;
    wire w558;
    wire w559;
    wire w560;
    wire w561;
    wire w562;
    wire w563;
    wire w564;
    wire w565;
    wire w566;
    assign out2[0] = w497;
    assign out2[1] = w498;
    assign out2[2] = w499;
    assign out2[3] = w500;
    assign out2[4] = w501;
    assign out2[5] = w502;
    assign out2[6] = w503;
    assign out2[7] = w504;
    assign out2[8] = w505;
    assign out2[9] = w506;
    assign out2[10] = w507;
    assign out2[11] = w508;
    assign out2[12] = w509;
    assign out2[13] = w510;
    assign out2[14] = w511;
    assign out2[15] = w512;
    assign out2[16] = w513;
    assign out2[17] = w514;
    assign out2[18] = w515;
    assign out2[19] = w516;
    assign out2[20] = w517;
    assign out2[21] = w518;
    assign out2[22] = w519;
    assign out2[23] = w520;
    assign out2[24] = w521;
    assign out2[25] = w522;
    assign out2[26] = w523;
    assign out2[27] = w524;
    assign out2[28] = w525;
    assign out2[29] = w526;
    assign out2[30] = w527;
    assign out2[31] = w528;
    assign out2[32] = w529;
    assign out2[33] = w530;
    assign out2[34] = w531;
    assign out2[35] = w532;
    assign out2[36] = w533;
    assign out2[37] = w534;
    assign out2[38] = w535;
    assign out2[39] = w536;
    assign out2[40] = w537;
    assign out2[41] = w538;
    assign out2[42] = w539;
    assign out2[43] = w540;
    assign out2[44] = w541;
    assign out2[45] = w542;
    assign out2[46] = w543;
    assign out2[47] = w544;
    assign out2[48] = w545;
    assign out2[49] = w546;
    assign out2[50] = w547;
    assign out2[51] = w548;
    assign out2[52] = w549;
    assign out2[53] = w550;
    assign out2[54] = w551;
    assign out2[55] = w552;
    assign out2[56] = w553;
    assign out2[57] = w554;
    assign out2[58] = w555;
    assign out2[59] = w556;
    assign out2[60] = w557;
    assign out2[61] = w558;
    assign out2[62] = w559;
    assign out2[63] = w560;
    assign out2[64] = w561;
    assign out2[65] = w562;
    assign out2[66] = w563;
    assign out2[67] = w564;
    assign out2[68] = w565;
    assign out2[69] = w566;
    wire w357;
    wire w358;
    wire w359;
    wire w360;
    wire w361;
    wire w362;
    wire w363;
    wire w364;
    wire w365;
    wire w366;
    wire w367;
    wire w368;
    wire w369;
    wire w370;
    wire w371;
    wire w372;
    wire w373;
    wire w374;
    wire w375;
    wire w376;
    wire w377;
    wire w378;
    wire w379;
    wire w380;
    wire w381;
    wire w382;
    wire w383;
    wire w384;
    wire w385;
    wire w386;
    wire w387;
    wire w388;
    wire w389;
    wire w390;
    wire w391;
    wire w392;
    wire w393;
    wire w394;
    wire w395;
    wire w396;
    wire w397;
    wire w398;
    wire w399;
    wire w400;
    wire w401;
    wire w402;
    wire w403;
    wire w404;
    wire w405;
    wire w406;
    wire w407;
    wire w408;
    wire w409;
    wire w410;
    wire w411;
    wire w412;
    wire w413;
    wire w414;
    wire w415;
    wire w416;
    wire w417;
    wire w418;
    wire w419;
    wire w420;
    wire w421;
    wire w422;
    wire w423;
    wire w424;
    wire w425;
    wire w426;
    assign out3[0] = w357;
    assign out3[1] = w358;
    assign out3[2] = w359;
    assign out3[3] = w360;
    assign out3[4] = w361;
    assign out3[5] = w362;
    assign out3[6] = w363;
    assign out3[7] = w364;
    assign out3[8] = w365;
    assign out3[9] = w366;
    assign out3[10] = w367;
    assign out3[11] = w368;
    assign out3[12] = w369;
    assign out3[13] = w370;
    assign out3[14] = w371;
    assign out3[15] = w372;
    assign out3[16] = w373;
    assign out3[17] = w374;
    assign out3[18] = w375;
    assign out3[19] = w376;
    assign out3[20] = w377;
    assign out3[21] = w378;
    assign out3[22] = w379;
    assign out3[23] = w380;
    assign out3[24] = w381;
    assign out3[25] = w382;
    assign out3[26] = w383;
    assign out3[27] = w384;
    assign out3[28] = w385;
    assign out3[29] = w386;
    assign out3[30] = w387;
    assign out3[31] = w388;
    assign out3[32] = w389;
    assign out3[33] = w390;
    assign out3[34] = w391;
    assign out3[35] = w392;
    assign out3[36] = w393;
    assign out3[37] = w394;
    assign out3[38] = w395;
    assign out3[39] = w396;
    assign out3[40] = w397;
    assign out3[41] = w398;
    assign out3[42] = w399;
    assign out3[43] = w400;
    assign out3[44] = w401;
    assign out3[45] = w402;
    assign out3[46] = w403;
    assign out3[47] = w404;
    assign out3[48] = w405;
    assign out3[49] = w406;
    assign out3[50] = w407;
    assign out3[51] = w408;
    assign out3[52] = w409;
    assign out3[53] = w410;
    assign out3[54] = w411;
    assign out3[55] = w412;
    assign out3[56] = w413;
    assign out3[57] = w414;
    assign out3[58] = w415;
    assign out3[59] = w416;
    assign out3[60] = w417;
    assign out3[61] = w418;
    assign out3[62] = w419;
    assign out3[63] = w420;
    assign out3[64] = w421;
    assign out3[65] = w422;
    assign out3[66] = w423;
    assign out3[67] = w424;
    assign out3[68] = w425;
    assign out3[69] = w426;
    wire w853;
    wire w854;
    wire w855;
    wire w856;
    wire w857;
    wire w858;
    wire w859;
    wire w860;
    wire w861;
    wire w862;
    wire w863;
    wire w864;
    wire w865;
    wire w866;
    wire w867;
    wire w868;
    wire w869;
    wire w870;
    wire w871;
    wire w872;
    wire w873;
    wire w874;
    wire w875;
    wire w876;
    wire w877;
    wire w878;
    wire w879;
    wire w880;
    wire w881;
    wire w882;
    wire w883;
    wire w884;
    wire w885;
    wire w886;
    wire w887;
    wire w888;
    wire w889;
    wire w890;
    wire w891;
    wire w892;
    wire w893;
    wire w894;
    wire w895;
    wire w896;
    wire w897;
    wire w898;
    wire w899;
    wire w900;
    wire w901;
    wire w902;
    wire w903;
    wire w904;
    wire w905;
    wire w906;
    wire w907;
    wire w908;
    wire w909;
    wire w910;
    wire w911;
    wire w912;
    wire w913;
    wire w914;
    wire w915;
    wire w916;
    wire w917;
    wire w918;
    wire w919;
    wire w920;
    wire w921;
    wire w922;
    assign out4[0] = w853;
    assign out4[1] = w854;
    assign out4[2] = w855;
    assign out4[3] = w856;
    assign out4[4] = w857;
    assign out4[5] = w858;
    assign out4[6] = w859;
    assign out4[7] = w860;
    assign out4[8] = w861;
    assign out4[9] = w862;
    assign out4[10] = w863;
    assign out4[11] = w864;
    assign out4[12] = w865;
    assign out4[13] = w866;
    assign out4[14] = w867;
    assign out4[15] = w868;
    assign out4[16] = w869;
    assign out4[17] = w870;
    assign out4[18] = w871;
    assign out4[19] = w872;
    assign out4[20] = w873;
    assign out4[21] = w874;
    assign out4[22] = w875;
    assign out4[23] = w876;
    assign out4[24] = w877;
    assign out4[25] = w878;
    assign out4[26] = w879;
    assign out4[27] = w880;
    assign out4[28] = w881;
    assign out4[29] = w882;
    assign out4[30] = w883;
    assign out4[31] = w884;
    assign out4[32] = w885;
    assign out4[33] = w886;
    assign out4[34] = w887;
    assign out4[35] = w888;
    assign out4[36] = w889;
    assign out4[37] = w890;
    assign out4[38] = w891;
    assign out4[39] = w892;
    assign out4[40] = w893;
    assign out4[41] = w894;
    assign out4[42] = w895;
    assign out4[43] = w896;
    assign out4[44] = w897;
    assign out4[45] = w898;
    assign out4[46] = w899;
    assign out4[47] = w900;
    assign out4[48] = w901;
    assign out4[49] = w902;
    assign out4[50] = w903;
    assign out4[51] = w904;
    assign out4[52] = w905;
    assign out4[53] = w906;
    assign out4[54] = w907;
    assign out4[55] = w908;
    assign out4[56] = w909;
    assign out4[57] = w910;
    assign out4[58] = w911;
    assign out4[59] = w912;
    assign out4[60] = w913;
    assign out4[61] = w914;
    assign out4[62] = w915;
    assign out4[63] = w916;
    assign out4[64] = w917;
    assign out4[65] = w918;
    assign out4[66] = w919;
    assign out4[67] = w920;
    assign out4[68] = w921;
    assign out4[69] = w922;
    wire w993;
    wire w994;
    wire w995;
    wire w996;
    wire w997;
    wire w998;
    wire w999;
    wire w1000;
    wire w1001;
    wire w1002;
    wire w1003;
    wire w1004;
    wire w1005;
    wire w1006;
    wire w1007;
    wire w1008;
    wire w1009;
    wire w1010;
    wire w1011;
    wire w1012;
    wire w1013;
    wire w1014;
    wire w1015;
    wire w1016;
    wire w1017;
    wire w1018;
    wire w1019;
    wire w1020;
    wire w1021;
    wire w1022;
    wire w1023;
    wire w1024;
    wire w1025;
    wire w1026;
    wire w1027;
    wire w1028;
    wire w1029;
    wire w1030;
    wire w1031;
    wire w1032;
    wire w1033;
    wire w1034;
    wire w1035;
    wire w1036;
    wire w1037;
    wire w1038;
    wire w1039;
    wire w1040;
    wire w1041;
    wire w1042;
    wire w1043;
    wire w1044;
    wire w1045;
    wire w1046;
    wire w1047;
    wire w1048;
    wire w1049;
    wire w1050;
    wire w1051;
    wire w1052;
    wire w1053;
    wire w1054;
    wire w1055;
    wire w1056;
    wire w1057;
    wire w1058;
    wire w1059;
    wire w1060;
    wire w1061;
    wire w1062;
    assign out5[0] = w993;
    assign out5[1] = w994;
    assign out5[2] = w995;
    assign out5[3] = w996;
    assign out5[4] = w997;
    assign out5[5] = w998;
    assign out5[6] = w999;
    assign out5[7] = w1000;
    assign out5[8] = w1001;
    assign out5[9] = w1002;
    assign out5[10] = w1003;
    assign out5[11] = w1004;
    assign out5[12] = w1005;
    assign out5[13] = w1006;
    assign out5[14] = w1007;
    assign out5[15] = w1008;
    assign out5[16] = w1009;
    assign out5[17] = w1010;
    assign out5[18] = w1011;
    assign out5[19] = w1012;
    assign out5[20] = w1013;
    assign out5[21] = w1014;
    assign out5[22] = w1015;
    assign out5[23] = w1016;
    assign out5[24] = w1017;
    assign out5[25] = w1018;
    assign out5[26] = w1019;
    assign out5[27] = w1020;
    assign out5[28] = w1021;
    assign out5[29] = w1022;
    assign out5[30] = w1023;
    assign out5[31] = w1024;
    assign out5[32] = w1025;
    assign out5[33] = w1026;
    assign out5[34] = w1027;
    assign out5[35] = w1028;
    assign out5[36] = w1029;
    assign out5[37] = w1030;
    assign out5[38] = w1031;
    assign out5[39] = w1032;
    assign out5[40] = w1033;
    assign out5[41] = w1034;
    assign out5[42] = w1035;
    assign out5[43] = w1036;
    assign out5[44] = w1037;
    assign out5[45] = w1038;
    assign out5[46] = w1039;
    assign out5[47] = w1040;
    assign out5[48] = w1041;
    assign out5[49] = w1042;
    assign out5[50] = w1043;
    assign out5[51] = w1044;
    assign out5[52] = w1045;
    assign out5[53] = w1046;
    assign out5[54] = w1047;
    assign out5[55] = w1048;
    assign out5[56] = w1049;
    assign out5[57] = w1050;
    assign out5[58] = w1051;
    assign out5[59] = w1052;
    assign out5[60] = w1053;
    assign out5[61] = w1054;
    assign out5[62] = w1055;
    assign out5[63] = w1056;
    assign out5[64] = w1057;
    assign out5[65] = w1058;
    assign out5[66] = w1059;
    assign out5[67] = w1060;
    assign out5[68] = w1061;
    assign out5[69] = w1062;
    wire w1063;
    wire w1064;
    wire w1065;
    wire w1066;
    wire w1067;
    wire w1068;
    wire w1069;
    wire w1070;
    wire w1071;
    wire w1072;
    wire w1073;
    wire w1074;
    wire w1075;
    wire w1076;
    wire w1077;
    wire w1078;
    wire w1079;
    wire w1080;
    wire w1081;
    wire w1082;
    wire w1083;
    wire w1084;
    wire w1085;
    wire w1086;
    wire w1087;
    wire w1088;
    wire w1089;
    wire w1090;
    wire w1091;
    wire w1092;
    wire w1093;
    wire w1094;
    wire w1095;
    wire w1096;
    wire w1097;
    wire w1098;
    wire w1099;
    wire w1100;
    wire w1101;
    wire w1102;
    wire w1103;
    wire w1104;
    wire w1105;
    wire w1106;
    wire w1107;
    wire w1108;
    wire w1109;
    wire w1110;
    wire w1111;
    wire w1112;
    wire w1113;
    wire w1114;
    wire w1115;
    wire w1116;
    wire w1117;
    wire w1118;
    wire w1119;
    wire w1120;
    wire w1121;
    wire w1122;
    wire w1123;
    wire w1124;
    wire w1125;
    wire w1126;
    wire w1127;
    wire w1128;
    wire w1129;
    wire w1130;
    wire w1131;
    wire w1132;
    assign out6[0] = w1063;
    assign out6[1] = w1064;
    assign out6[2] = w1065;
    assign out6[3] = w1066;
    assign out6[4] = w1067;
    assign out6[5] = w1068;
    assign out6[6] = w1069;
    assign out6[7] = w1070;
    assign out6[8] = w1071;
    assign out6[9] = w1072;
    assign out6[10] = w1073;
    assign out6[11] = w1074;
    assign out6[12] = w1075;
    assign out6[13] = w1076;
    assign out6[14] = w1077;
    assign out6[15] = w1078;
    assign out6[16] = w1079;
    assign out6[17] = w1080;
    assign out6[18] = w1081;
    assign out6[19] = w1082;
    assign out6[20] = w1083;
    assign out6[21] = w1084;
    assign out6[22] = w1085;
    assign out6[23] = w1086;
    assign out6[24] = w1087;
    assign out6[25] = w1088;
    assign out6[26] = w1089;
    assign out6[27] = w1090;
    assign out6[28] = w1091;
    assign out6[29] = w1092;
    assign out6[30] = w1093;
    assign out6[31] = w1094;
    assign out6[32] = w1095;
    assign out6[33] = w1096;
    assign out6[34] = w1097;
    assign out6[35] = w1098;
    assign out6[36] = w1099;
    assign out6[37] = w1100;
    assign out6[38] = w1101;
    assign out6[39] = w1102;
    assign out6[40] = w1103;
    assign out6[41] = w1104;
    assign out6[42] = w1105;
    assign out6[43] = w1106;
    assign out6[44] = w1107;
    assign out6[45] = w1108;
    assign out6[46] = w1109;
    assign out6[47] = w1110;
    assign out6[48] = w1111;
    assign out6[49] = w1112;
    assign out6[50] = w1113;
    assign out6[51] = w1114;
    assign out6[52] = w1115;
    assign out6[53] = w1116;
    assign out6[54] = w1117;
    assign out6[55] = w1118;
    assign out6[56] = w1119;
    assign out6[57] = w1120;
    assign out6[58] = w1121;
    assign out6[59] = w1122;
    assign out6[60] = w1123;
    assign out6[61] = w1124;
    assign out6[62] = w1125;
    assign out6[63] = w1126;
    assign out6[64] = w1127;
    assign out6[65] = w1128;
    assign out6[66] = w1129;
    assign out6[67] = w1130;
    assign out6[68] = w1131;
    assign out6[69] = w1132;
    wire w923;
    wire w924;
    wire w925;
    wire w926;
    wire w927;
    wire w928;
    wire w929;
    wire w930;
    wire w931;
    wire w932;
    wire w933;
    wire w934;
    wire w935;
    wire w936;
    wire w937;
    wire w938;
    wire w939;
    wire w940;
    wire w941;
    wire w942;
    wire w943;
    wire w944;
    wire w945;
    wire w946;
    wire w947;
    wire w948;
    wire w949;
    wire w950;
    wire w951;
    wire w952;
    wire w953;
    wire w954;
    wire w955;
    wire w956;
    wire w957;
    wire w958;
    wire w959;
    wire w960;
    wire w961;
    wire w962;
    wire w963;
    wire w964;
    wire w965;
    wire w966;
    wire w967;
    wire w968;
    wire w969;
    wire w970;
    wire w971;
    wire w972;
    wire w973;
    wire w974;
    wire w975;
    wire w976;
    wire w977;
    wire w978;
    wire w979;
    wire w980;
    wire w981;
    wire w982;
    wire w983;
    wire w984;
    wire w985;
    wire w986;
    wire w987;
    wire w988;
    wire w989;
    wire w990;
    wire w991;
    wire w992;
    assign out7[0] = w923;
    assign out7[1] = w924;
    assign out7[2] = w925;
    assign out7[3] = w926;
    assign out7[4] = w927;
    assign out7[5] = w928;
    assign out7[6] = w929;
    assign out7[7] = w930;
    assign out7[8] = w931;
    assign out7[9] = w932;
    assign out7[10] = w933;
    assign out7[11] = w934;
    assign out7[12] = w935;
    assign out7[13] = w936;
    assign out7[14] = w937;
    assign out7[15] = w938;
    assign out7[16] = w939;
    assign out7[17] = w940;
    assign out7[18] = w941;
    assign out7[19] = w942;
    assign out7[20] = w943;
    assign out7[21] = w944;
    assign out7[22] = w945;
    assign out7[23] = w946;
    assign out7[24] = w947;
    assign out7[25] = w948;
    assign out7[26] = w949;
    assign out7[27] = w950;
    assign out7[28] = w951;
    assign out7[29] = w952;
    assign out7[30] = w953;
    assign out7[31] = w954;
    assign out7[32] = w955;
    assign out7[33] = w956;
    assign out7[34] = w957;
    assign out7[35] = w958;
    assign out7[36] = w959;
    assign out7[37] = w960;
    assign out7[38] = w961;
    assign out7[39] = w962;
    assign out7[40] = w963;
    assign out7[41] = w964;
    assign out7[42] = w965;
    assign out7[43] = w966;
    assign out7[44] = w967;
    assign out7[45] = w968;
    assign out7[46] = w969;
    assign out7[47] = w970;
    assign out7[48] = w971;
    assign out7[49] = w972;
    assign out7[50] = w973;
    assign out7[51] = w974;
    assign out7[52] = w975;
    assign out7[53] = w976;
    assign out7[54] = w977;
    assign out7[55] = w978;
    assign out7[56] = w979;
    assign out7[57] = w980;
    assign out7[58] = w981;
    assign out7[59] = w982;
    assign out7[60] = w983;
    assign out7[61] = w984;
    assign out7[62] = w985;
    assign out7[63] = w986;
    assign out7[64] = w987;
    assign out7[65] = w988;
    assign out7[66] = w989;
    assign out7[67] = w990;
    assign out7[68] = w991;
    assign out7[69] = w992;
    wire w1419;
    wire w1420;
    wire w1421;
    wire w1422;
    wire w1423;
    wire w1424;
    wire w1425;
    wire w1426;
    wire w1427;
    wire w1428;
    wire w1429;
    wire w1430;
    wire w1431;
    wire w1432;
    wire w1433;
    wire w1434;
    wire w1435;
    wire w1436;
    wire w1437;
    wire w1438;
    wire w1439;
    wire w1440;
    wire w1441;
    wire w1442;
    wire w1443;
    wire w1444;
    wire w1445;
    wire w1446;
    wire w1447;
    wire w1448;
    wire w1449;
    wire w1450;
    wire w1451;
    wire w1452;
    wire w1453;
    wire w1454;
    wire w1455;
    wire w1456;
    wire w1457;
    wire w1458;
    wire w1459;
    wire w1460;
    wire w1461;
    wire w1462;
    wire w1463;
    wire w1464;
    wire w1465;
    wire w1466;
    wire w1467;
    wire w1468;
    wire w1469;
    wire w1470;
    wire w1471;
    wire w1472;
    wire w1473;
    wire w1474;
    wire w1475;
    wire w1476;
    wire w1477;
    wire w1478;
    wire w1479;
    wire w1480;
    wire w1481;
    wire w1482;
    wire w1483;
    wire w1484;
    wire w1485;
    wire w1486;
    wire w1487;
    wire w1488;
    assign out8[0] = w1419;
    assign out8[1] = w1420;
    assign out8[2] = w1421;
    assign out8[3] = w1422;
    assign out8[4] = w1423;
    assign out8[5] = w1424;
    assign out8[6] = w1425;
    assign out8[7] = w1426;
    assign out8[8] = w1427;
    assign out8[9] = w1428;
    assign out8[10] = w1429;
    assign out8[11] = w1430;
    assign out8[12] = w1431;
    assign out8[13] = w1432;
    assign out8[14] = w1433;
    assign out8[15] = w1434;
    assign out8[16] = w1435;
    assign out8[17] = w1436;
    assign out8[18] = w1437;
    assign out8[19] = w1438;
    assign out8[20] = w1439;
    assign out8[21] = w1440;
    assign out8[22] = w1441;
    assign out8[23] = w1442;
    assign out8[24] = w1443;
    assign out8[25] = w1444;
    assign out8[26] = w1445;
    assign out8[27] = w1446;
    assign out8[28] = w1447;
    assign out8[29] = w1448;
    assign out8[30] = w1449;
    assign out8[31] = w1450;
    assign out8[32] = w1451;
    assign out8[33] = w1452;
    assign out8[34] = w1453;
    assign out8[35] = w1454;
    assign out8[36] = w1455;
    assign out8[37] = w1456;
    assign out8[38] = w1457;
    assign out8[39] = w1458;
    assign out8[40] = w1459;
    assign out8[41] = w1460;
    assign out8[42] = w1461;
    assign out8[43] = w1462;
    assign out8[44] = w1463;
    assign out8[45] = w1464;
    assign out8[46] = w1465;
    assign out8[47] = w1466;
    assign out8[48] = w1467;
    assign out8[49] = w1468;
    assign out8[50] = w1469;
    assign out8[51] = w1470;
    assign out8[52] = w1471;
    assign out8[53] = w1472;
    assign out8[54] = w1473;
    assign out8[55] = w1474;
    assign out8[56] = w1475;
    assign out8[57] = w1476;
    assign out8[58] = w1477;
    assign out8[59] = w1478;
    assign out8[60] = w1479;
    assign out8[61] = w1480;
    assign out8[62] = w1481;
    assign out8[63] = w1482;
    assign out8[64] = w1483;
    assign out8[65] = w1484;
    assign out8[66] = w1485;
    assign out8[67] = w1486;
    assign out8[68] = w1487;
    assign out8[69] = w1488;
    wire w1559;
    wire w1560;
    wire w1561;
    wire w1562;
    wire w1563;
    wire w1564;
    wire w1565;
    wire w1566;
    wire w1567;
    wire w1568;
    wire w1569;
    wire w1570;
    wire w1571;
    wire w1572;
    wire w1573;
    wire w1574;
    wire w1575;
    wire w1576;
    wire w1577;
    wire w1578;
    wire w1579;
    wire w1580;
    wire w1581;
    wire w1582;
    wire w1583;
    wire w1584;
    wire w1585;
    wire w1586;
    wire w1587;
    wire w1588;
    wire w1589;
    wire w1590;
    wire w1591;
    wire w1592;
    wire w1593;
    wire w1594;
    wire w1595;
    wire w1596;
    wire w1597;
    wire w1598;
    wire w1599;
    wire w1600;
    wire w1601;
    wire w1602;
    wire w1603;
    wire w1604;
    wire w1605;
    wire w1606;
    wire w1607;
    wire w1608;
    wire w1609;
    wire w1610;
    wire w1611;
    wire w1612;
    wire w1613;
    wire w1614;
    wire w1615;
    wire w1616;
    wire w1617;
    wire w1618;
    wire w1619;
    wire w1620;
    wire w1621;
    wire w1622;
    wire w1623;
    wire w1624;
    wire w1625;
    wire w1626;
    wire w1627;
    wire w1628;
    assign out9[0] = w1559;
    assign out9[1] = w1560;
    assign out9[2] = w1561;
    assign out9[3] = w1562;
    assign out9[4] = w1563;
    assign out9[5] = w1564;
    assign out9[6] = w1565;
    assign out9[7] = w1566;
    assign out9[8] = w1567;
    assign out9[9] = w1568;
    assign out9[10] = w1569;
    assign out9[11] = w1570;
    assign out9[12] = w1571;
    assign out9[13] = w1572;
    assign out9[14] = w1573;
    assign out9[15] = w1574;
    assign out9[16] = w1575;
    assign out9[17] = w1576;
    assign out9[18] = w1577;
    assign out9[19] = w1578;
    assign out9[20] = w1579;
    assign out9[21] = w1580;
    assign out9[22] = w1581;
    assign out9[23] = w1582;
    assign out9[24] = w1583;
    assign out9[25] = w1584;
    assign out9[26] = w1585;
    assign out9[27] = w1586;
    assign out9[28] = w1587;
    assign out9[29] = w1588;
    assign out9[30] = w1589;
    assign out9[31] = w1590;
    assign out9[32] = w1591;
    assign out9[33] = w1592;
    assign out9[34] = w1593;
    assign out9[35] = w1594;
    assign out9[36] = w1595;
    assign out9[37] = w1596;
    assign out9[38] = w1597;
    assign out9[39] = w1598;
    assign out9[40] = w1599;
    assign out9[41] = w1600;
    assign out9[42] = w1601;
    assign out9[43] = w1602;
    assign out9[44] = w1603;
    assign out9[45] = w1604;
    assign out9[46] = w1605;
    assign out9[47] = w1606;
    assign out9[48] = w1607;
    assign out9[49] = w1608;
    assign out9[50] = w1609;
    assign out9[51] = w1610;
    assign out9[52] = w1611;
    assign out9[53] = w1612;
    assign out9[54] = w1613;
    assign out9[55] = w1614;
    assign out9[56] = w1615;
    assign out9[57] = w1616;
    assign out9[58] = w1617;
    assign out9[59] = w1618;
    assign out9[60] = w1619;
    assign out9[61] = w1620;
    assign out9[62] = w1621;
    assign out9[63] = w1622;
    assign out9[64] = w1623;
    assign out9[65] = w1624;
    assign out9[66] = w1625;
    assign out9[67] = w1626;
    assign out9[68] = w1627;
    assign out9[69] = w1628;
    wire w1629;
    wire w1630;
    wire w1631;
    wire w1632;
    wire w1633;
    wire w1634;
    wire w1635;
    wire w1636;
    wire w1637;
    wire w1638;
    wire w1639;
    wire w1640;
    wire w1641;
    wire w1642;
    wire w1643;
    wire w1644;
    wire w1645;
    wire w1646;
    wire w1647;
    wire w1648;
    wire w1649;
    wire w1650;
    wire w1651;
    wire w1652;
    wire w1653;
    wire w1654;
    wire w1655;
    wire w1656;
    wire w1657;
    wire w1658;
    wire w1659;
    wire w1660;
    wire w1661;
    wire w1662;
    wire w1663;
    wire w1664;
    wire w1665;
    wire w1666;
    wire w1667;
    wire w1668;
    wire w1669;
    wire w1670;
    wire w1671;
    wire w1672;
    wire w1673;
    wire w1674;
    wire w1675;
    wire w1676;
    wire w1677;
    wire w1678;
    wire w1679;
    wire w1680;
    wire w1681;
    wire w1682;
    wire w1683;
    wire w1684;
    wire w1685;
    wire w1686;
    wire w1687;
    wire w1688;
    wire w1689;
    wire w1690;
    wire w1691;
    wire w1692;
    wire w1693;
    wire w1694;
    wire w1695;
    wire w1696;
    wire w1697;
    wire w1698;
    assign out10[0] = w1629;
    assign out10[1] = w1630;
    assign out10[2] = w1631;
    assign out10[3] = w1632;
    assign out10[4] = w1633;
    assign out10[5] = w1634;
    assign out10[6] = w1635;
    assign out10[7] = w1636;
    assign out10[8] = w1637;
    assign out10[9] = w1638;
    assign out10[10] = w1639;
    assign out10[11] = w1640;
    assign out10[12] = w1641;
    assign out10[13] = w1642;
    assign out10[14] = w1643;
    assign out10[15] = w1644;
    assign out10[16] = w1645;
    assign out10[17] = w1646;
    assign out10[18] = w1647;
    assign out10[19] = w1648;
    assign out10[20] = w1649;
    assign out10[21] = w1650;
    assign out10[22] = w1651;
    assign out10[23] = w1652;
    assign out10[24] = w1653;
    assign out10[25] = w1654;
    assign out10[26] = w1655;
    assign out10[27] = w1656;
    assign out10[28] = w1657;
    assign out10[29] = w1658;
    assign out10[30] = w1659;
    assign out10[31] = w1660;
    assign out10[32] = w1661;
    assign out10[33] = w1662;
    assign out10[34] = w1663;
    assign out10[35] = w1664;
    assign out10[36] = w1665;
    assign out10[37] = w1666;
    assign out10[38] = w1667;
    assign out10[39] = w1668;
    assign out10[40] = w1669;
    assign out10[41] = w1670;
    assign out10[42] = w1671;
    assign out10[43] = w1672;
    assign out10[44] = w1673;
    assign out10[45] = w1674;
    assign out10[46] = w1675;
    assign out10[47] = w1676;
    assign out10[48] = w1677;
    assign out10[49] = w1678;
    assign out10[50] = w1679;
    assign out10[51] = w1680;
    assign out10[52] = w1681;
    assign out10[53] = w1682;
    assign out10[54] = w1683;
    assign out10[55] = w1684;
    assign out10[56] = w1685;
    assign out10[57] = w1686;
    assign out10[58] = w1687;
    assign out10[59] = w1688;
    assign out10[60] = w1689;
    assign out10[61] = w1690;
    assign out10[62] = w1691;
    assign out10[63] = w1692;
    assign out10[64] = w1693;
    assign out10[65] = w1694;
    assign out10[66] = w1695;
    assign out10[67] = w1696;
    assign out10[68] = w1697;
    assign out10[69] = w1698;
    wire w1489;
    wire w1490;
    wire w1491;
    wire w1492;
    wire w1493;
    wire w1494;
    wire w1495;
    wire w1496;
    wire w1497;
    wire w1498;
    wire w1499;
    wire w1500;
    wire w1501;
    wire w1502;
    wire w1503;
    wire w1504;
    wire w1505;
    wire w1506;
    wire w1507;
    wire w1508;
    wire w1509;
    wire w1510;
    wire w1511;
    wire w1512;
    wire w1513;
    wire w1514;
    wire w1515;
    wire w1516;
    wire w1517;
    wire w1518;
    wire w1519;
    wire w1520;
    wire w1521;
    wire w1522;
    wire w1523;
    wire w1524;
    wire w1525;
    wire w1526;
    wire w1527;
    wire w1528;
    wire w1529;
    wire w1530;
    wire w1531;
    wire w1532;
    wire w1533;
    wire w1534;
    wire w1535;
    wire w1536;
    wire w1537;
    wire w1538;
    wire w1539;
    wire w1540;
    wire w1541;
    wire w1542;
    wire w1543;
    wire w1544;
    wire w1545;
    wire w1546;
    wire w1547;
    wire w1548;
    wire w1549;
    wire w1550;
    wire w1551;
    wire w1552;
    wire w1553;
    wire w1554;
    wire w1555;
    wire w1556;
    wire w1557;
    wire w1558;
    assign out11[0] = w1489;
    assign out11[1] = w1490;
    assign out11[2] = w1491;
    assign out11[3] = w1492;
    assign out11[4] = w1493;
    assign out11[5] = w1494;
    assign out11[6] = w1495;
    assign out11[7] = w1496;
    assign out11[8] = w1497;
    assign out11[9] = w1498;
    assign out11[10] = w1499;
    assign out11[11] = w1500;
    assign out11[12] = w1501;
    assign out11[13] = w1502;
    assign out11[14] = w1503;
    assign out11[15] = w1504;
    assign out11[16] = w1505;
    assign out11[17] = w1506;
    assign out11[18] = w1507;
    assign out11[19] = w1508;
    assign out11[20] = w1509;
    assign out11[21] = w1510;
    assign out11[22] = w1511;
    assign out11[23] = w1512;
    assign out11[24] = w1513;
    assign out11[25] = w1514;
    assign out11[26] = w1515;
    assign out11[27] = w1516;
    assign out11[28] = w1517;
    assign out11[29] = w1518;
    assign out11[30] = w1519;
    assign out11[31] = w1520;
    assign out11[32] = w1521;
    assign out11[33] = w1522;
    assign out11[34] = w1523;
    assign out11[35] = w1524;
    assign out11[36] = w1525;
    assign out11[37] = w1526;
    assign out11[38] = w1527;
    assign out11[39] = w1528;
    assign out11[40] = w1529;
    assign out11[41] = w1530;
    assign out11[42] = w1531;
    assign out11[43] = w1532;
    assign out11[44] = w1533;
    assign out11[45] = w1534;
    assign out11[46] = w1535;
    assign out11[47] = w1536;
    assign out11[48] = w1537;
    assign out11[49] = w1538;
    assign out11[50] = w1539;
    assign out11[51] = w1540;
    assign out11[52] = w1541;
    assign out11[53] = w1542;
    assign out11[54] = w1543;
    assign out11[55] = w1544;
    assign out11[56] = w1545;
    assign out11[57] = w1546;
    assign out11[58] = w1547;
    assign out11[59] = w1548;
    assign out11[60] = w1549;
    assign out11[61] = w1550;
    assign out11[62] = w1551;
    assign out11[63] = w1552;
    assign out11[64] = w1553;
    assign out11[65] = w1554;
    assign out11[66] = w1555;
    assign out11[67] = w1556;
    assign out11[68] = w1557;
    assign out11[69] = w1558;
    wire w1985;
    wire w1986;
    wire w1987;
    wire w1988;
    wire w1989;
    wire w1990;
    wire w1991;
    wire w1992;
    wire w1993;
    wire w1994;
    wire w1995;
    wire w1996;
    wire w1997;
    wire w1998;
    wire w1999;
    wire w2000;
    wire w2001;
    wire w2002;
    wire w2003;
    wire w2004;
    wire w2005;
    wire w2006;
    wire w2007;
    wire w2008;
    wire w2009;
    wire w2010;
    wire w2011;
    wire w2012;
    wire w2013;
    wire w2014;
    wire w2015;
    wire w2016;
    wire w2017;
    wire w2018;
    wire w2019;
    wire w2020;
    wire w2021;
    wire w2022;
    wire w2023;
    wire w2024;
    wire w2025;
    wire w2026;
    wire w2027;
    wire w2028;
    wire w2029;
    wire w2030;
    wire w2031;
    wire w2032;
    wire w2033;
    wire w2034;
    wire w2035;
    wire w2036;
    wire w2037;
    wire w2038;
    wire w2039;
    wire w2040;
    wire w2041;
    wire w2042;
    wire w2043;
    wire w2044;
    wire w2045;
    wire w2046;
    wire w2047;
    wire w2048;
    wire w2049;
    wire w2050;
    wire w2051;
    wire w2052;
    wire w2053;
    wire w2054;
    assign out12[0] = w1985;
    assign out12[1] = w1986;
    assign out12[2] = w1987;
    assign out12[3] = w1988;
    assign out12[4] = w1989;
    assign out12[5] = w1990;
    assign out12[6] = w1991;
    assign out12[7] = w1992;
    assign out12[8] = w1993;
    assign out12[9] = w1994;
    assign out12[10] = w1995;
    assign out12[11] = w1996;
    assign out12[12] = w1997;
    assign out12[13] = w1998;
    assign out12[14] = w1999;
    assign out12[15] = w2000;
    assign out12[16] = w2001;
    assign out12[17] = w2002;
    assign out12[18] = w2003;
    assign out12[19] = w2004;
    assign out12[20] = w2005;
    assign out12[21] = w2006;
    assign out12[22] = w2007;
    assign out12[23] = w2008;
    assign out12[24] = w2009;
    assign out12[25] = w2010;
    assign out12[26] = w2011;
    assign out12[27] = w2012;
    assign out12[28] = w2013;
    assign out12[29] = w2014;
    assign out12[30] = w2015;
    assign out12[31] = w2016;
    assign out12[32] = w2017;
    assign out12[33] = w2018;
    assign out12[34] = w2019;
    assign out12[35] = w2020;
    assign out12[36] = w2021;
    assign out12[37] = w2022;
    assign out12[38] = w2023;
    assign out12[39] = w2024;
    assign out12[40] = w2025;
    assign out12[41] = w2026;
    assign out12[42] = w2027;
    assign out12[43] = w2028;
    assign out12[44] = w2029;
    assign out12[45] = w2030;
    assign out12[46] = w2031;
    assign out12[47] = w2032;
    assign out12[48] = w2033;
    assign out12[49] = w2034;
    assign out12[50] = w2035;
    assign out12[51] = w2036;
    assign out12[52] = w2037;
    assign out12[53] = w2038;
    assign out12[54] = w2039;
    assign out12[55] = w2040;
    assign out12[56] = w2041;
    assign out12[57] = w2042;
    assign out12[58] = w2043;
    assign out12[59] = w2044;
    assign out12[60] = w2045;
    assign out12[61] = w2046;
    assign out12[62] = w2047;
    assign out12[63] = w2048;
    assign out12[64] = w2049;
    assign out12[65] = w2050;
    assign out12[66] = w2051;
    assign out12[67] = w2052;
    assign out12[68] = w2053;
    assign out12[69] = w2054;
    wire w2125;
    wire w2126;
    wire w2127;
    wire w2128;
    wire w2129;
    wire w2130;
    wire w2131;
    wire w2132;
    wire w2133;
    wire w2134;
    wire w2135;
    wire w2136;
    wire w2137;
    wire w2138;
    wire w2139;
    wire w2140;
    wire w2141;
    wire w2142;
    wire w2143;
    wire w2144;
    wire w2145;
    wire w2146;
    wire w2147;
    wire w2148;
    wire w2149;
    wire w2150;
    wire w2151;
    wire w2152;
    wire w2153;
    wire w2154;
    wire w2155;
    wire w2156;
    wire w2157;
    wire w2158;
    wire w2159;
    wire w2160;
    wire w2161;
    wire w2162;
    wire w2163;
    wire w2164;
    wire w2165;
    wire w2166;
    wire w2167;
    wire w2168;
    wire w2169;
    wire w2170;
    wire w2171;
    wire w2172;
    wire w2173;
    wire w2174;
    wire w2175;
    wire w2176;
    wire w2177;
    wire w2178;
    wire w2179;
    wire w2180;
    wire w2181;
    wire w2182;
    wire w2183;
    wire w2184;
    wire w2185;
    wire w2186;
    wire w2187;
    wire w2188;
    wire w2189;
    wire w2190;
    wire w2191;
    wire w2192;
    wire w2193;
    wire w2194;
    assign out13[0] = w2125;
    assign out13[1] = w2126;
    assign out13[2] = w2127;
    assign out13[3] = w2128;
    assign out13[4] = w2129;
    assign out13[5] = w2130;
    assign out13[6] = w2131;
    assign out13[7] = w2132;
    assign out13[8] = w2133;
    assign out13[9] = w2134;
    assign out13[10] = w2135;
    assign out13[11] = w2136;
    assign out13[12] = w2137;
    assign out13[13] = w2138;
    assign out13[14] = w2139;
    assign out13[15] = w2140;
    assign out13[16] = w2141;
    assign out13[17] = w2142;
    assign out13[18] = w2143;
    assign out13[19] = w2144;
    assign out13[20] = w2145;
    assign out13[21] = w2146;
    assign out13[22] = w2147;
    assign out13[23] = w2148;
    assign out13[24] = w2149;
    assign out13[25] = w2150;
    assign out13[26] = w2151;
    assign out13[27] = w2152;
    assign out13[28] = w2153;
    assign out13[29] = w2154;
    assign out13[30] = w2155;
    assign out13[31] = w2156;
    assign out13[32] = w2157;
    assign out13[33] = w2158;
    assign out13[34] = w2159;
    assign out13[35] = w2160;
    assign out13[36] = w2161;
    assign out13[37] = w2162;
    assign out13[38] = w2163;
    assign out13[39] = w2164;
    assign out13[40] = w2165;
    assign out13[41] = w2166;
    assign out13[42] = w2167;
    assign out13[43] = w2168;
    assign out13[44] = w2169;
    assign out13[45] = w2170;
    assign out13[46] = w2171;
    assign out13[47] = w2172;
    assign out13[48] = w2173;
    assign out13[49] = w2174;
    assign out13[50] = w2175;
    assign out13[51] = w2176;
    assign out13[52] = w2177;
    assign out13[53] = w2178;
    assign out13[54] = w2179;
    assign out13[55] = w2180;
    assign out13[56] = w2181;
    assign out13[57] = w2182;
    assign out13[58] = w2183;
    assign out13[59] = w2184;
    assign out13[60] = w2185;
    assign out13[61] = w2186;
    assign out13[62] = w2187;
    assign out13[63] = w2188;
    assign out13[64] = w2189;
    assign out13[65] = w2190;
    assign out13[66] = w2191;
    assign out13[67] = w2192;
    assign out13[68] = w2193;
    assign out13[69] = w2194;
    wire w2195;
    wire w2196;
    wire w2197;
    wire w2198;
    wire w2199;
    wire w2200;
    wire w2201;
    wire w2202;
    wire w2203;
    wire w2204;
    wire w2205;
    wire w2206;
    wire w2207;
    wire w2208;
    wire w2209;
    wire w2210;
    wire w2211;
    wire w2212;
    wire w2213;
    wire w2214;
    wire w2215;
    wire w2216;
    wire w2217;
    wire w2218;
    wire w2219;
    wire w2220;
    wire w2221;
    wire w2222;
    wire w2223;
    wire w2224;
    wire w2225;
    wire w2226;
    wire w2227;
    wire w2228;
    wire w2229;
    wire w2230;
    wire w2231;
    wire w2232;
    wire w2233;
    wire w2234;
    wire w2235;
    wire w2236;
    wire w2237;
    wire w2238;
    wire w2239;
    wire w2240;
    wire w2241;
    wire w2242;
    wire w2243;
    wire w2244;
    wire w2245;
    wire w2246;
    wire w2247;
    wire w2248;
    wire w2249;
    wire w2250;
    wire w2251;
    wire w2252;
    wire w2253;
    wire w2254;
    wire w2255;
    wire w2256;
    wire w2257;
    wire w2258;
    wire w2259;
    wire w2260;
    wire w2261;
    wire w2262;
    wire w2263;
    wire w2264;
    assign out14[0] = w2195;
    assign out14[1] = w2196;
    assign out14[2] = w2197;
    assign out14[3] = w2198;
    assign out14[4] = w2199;
    assign out14[5] = w2200;
    assign out14[6] = w2201;
    assign out14[7] = w2202;
    assign out14[8] = w2203;
    assign out14[9] = w2204;
    assign out14[10] = w2205;
    assign out14[11] = w2206;
    assign out14[12] = w2207;
    assign out14[13] = w2208;
    assign out14[14] = w2209;
    assign out14[15] = w2210;
    assign out14[16] = w2211;
    assign out14[17] = w2212;
    assign out14[18] = w2213;
    assign out14[19] = w2214;
    assign out14[20] = w2215;
    assign out14[21] = w2216;
    assign out14[22] = w2217;
    assign out14[23] = w2218;
    assign out14[24] = w2219;
    assign out14[25] = w2220;
    assign out14[26] = w2221;
    assign out14[27] = w2222;
    assign out14[28] = w2223;
    assign out14[29] = w2224;
    assign out14[30] = w2225;
    assign out14[31] = w2226;
    assign out14[32] = w2227;
    assign out14[33] = w2228;
    assign out14[34] = w2229;
    assign out14[35] = w2230;
    assign out14[36] = w2231;
    assign out14[37] = w2232;
    assign out14[38] = w2233;
    assign out14[39] = w2234;
    assign out14[40] = w2235;
    assign out14[41] = w2236;
    assign out14[42] = w2237;
    assign out14[43] = w2238;
    assign out14[44] = w2239;
    assign out14[45] = w2240;
    assign out14[46] = w2241;
    assign out14[47] = w2242;
    assign out14[48] = w2243;
    assign out14[49] = w2244;
    assign out14[50] = w2245;
    assign out14[51] = w2246;
    assign out14[52] = w2247;
    assign out14[53] = w2248;
    assign out14[54] = w2249;
    assign out14[55] = w2250;
    assign out14[56] = w2251;
    assign out14[57] = w2252;
    assign out14[58] = w2253;
    assign out14[59] = w2254;
    assign out14[60] = w2255;
    assign out14[61] = w2256;
    assign out14[62] = w2257;
    assign out14[63] = w2258;
    assign out14[64] = w2259;
    assign out14[65] = w2260;
    assign out14[66] = w2261;
    assign out14[67] = w2262;
    assign out14[68] = w2263;
    assign out14[69] = w2264;
    wire w2055;
    wire w2056;
    wire w2057;
    wire w2058;
    wire w2059;
    wire w2060;
    wire w2061;
    wire w2062;
    wire w2063;
    wire w2064;
    wire w2065;
    wire w2066;
    wire w2067;
    wire w2068;
    wire w2069;
    wire w2070;
    wire w2071;
    wire w2072;
    wire w2073;
    wire w2074;
    wire w2075;
    wire w2076;
    wire w2077;
    wire w2078;
    wire w2079;
    wire w2080;
    wire w2081;
    wire w2082;
    wire w2083;
    wire w2084;
    wire w2085;
    wire w2086;
    wire w2087;
    wire w2088;
    wire w2089;
    wire w2090;
    wire w2091;
    wire w2092;
    wire w2093;
    wire w2094;
    wire w2095;
    wire w2096;
    wire w2097;
    wire w2098;
    wire w2099;
    wire w2100;
    wire w2101;
    wire w2102;
    wire w2103;
    wire w2104;
    wire w2105;
    wire w2106;
    wire w2107;
    wire w2108;
    wire w2109;
    wire w2110;
    wire w2111;
    wire w2112;
    wire w2113;
    wire w2114;
    wire w2115;
    wire w2116;
    wire w2117;
    wire w2118;
    wire w2119;
    wire w2120;
    wire w2121;
    wire w2122;
    wire w2123;
    wire w2124;
    assign out15[0] = w2055;
    assign out15[1] = w2056;
    assign out15[2] = w2057;
    assign out15[3] = w2058;
    assign out15[4] = w2059;
    assign out15[5] = w2060;
    assign out15[6] = w2061;
    assign out15[7] = w2062;
    assign out15[8] = w2063;
    assign out15[9] = w2064;
    assign out15[10] = w2065;
    assign out15[11] = w2066;
    assign out15[12] = w2067;
    assign out15[13] = w2068;
    assign out15[14] = w2069;
    assign out15[15] = w2070;
    assign out15[16] = w2071;
    assign out15[17] = w2072;
    assign out15[18] = w2073;
    assign out15[19] = w2074;
    assign out15[20] = w2075;
    assign out15[21] = w2076;
    assign out15[22] = w2077;
    assign out15[23] = w2078;
    assign out15[24] = w2079;
    assign out15[25] = w2080;
    assign out15[26] = w2081;
    assign out15[27] = w2082;
    assign out15[28] = w2083;
    assign out15[29] = w2084;
    assign out15[30] = w2085;
    assign out15[31] = w2086;
    assign out15[32] = w2087;
    assign out15[33] = w2088;
    assign out15[34] = w2089;
    assign out15[35] = w2090;
    assign out15[36] = w2091;
    assign out15[37] = w2092;
    assign out15[38] = w2093;
    assign out15[39] = w2094;
    assign out15[40] = w2095;
    assign out15[41] = w2096;
    assign out15[42] = w2097;
    assign out15[43] = w2098;
    assign out15[44] = w2099;
    assign out15[45] = w2100;
    assign out15[46] = w2101;
    assign out15[47] = w2102;
    assign out15[48] = w2103;
    assign out15[49] = w2104;
    assign out15[50] = w2105;
    assign out15[51] = w2106;
    assign out15[52] = w2107;
    assign out15[53] = w2108;
    assign out15[54] = w2109;
    assign out15[55] = w2110;
    assign out15[56] = w2111;
    assign out15[57] = w2112;
    assign out15[58] = w2113;
    assign out15[59] = w2114;
    assign out15[60] = w2115;
    assign out15[61] = w2116;
    assign out15[62] = w2117;
    assign out15[63] = w2118;
    assign out15[64] = w2119;
    assign out15[65] = w2120;
    assign out15[66] = w2121;
    assign out15[67] = w2122;
    assign out15[68] = w2123;
    assign out15[69] = w2124;
    wire w1699;
    xor xor0(w1699, x13_70, x14_70);
    wire w1;
    xor xor1(w1, x1_70, x2_70);
    wire w567;
    xor xor2(w567, x5_70, x6_70);
    wire w1133;
    xor xor3(w1133, x9_70, x10_70);
    wire w10, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w11, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w12, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w13, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w14, w140, w141, w142, w143, w144, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w3, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w4, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w5, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w6, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w7, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w8, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w9, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99;
    sw_m #(.SIZE(71)) sw4({w73,w72,w71,w70,w69,w68,w67,w66,w65,w64,w63,w62,w61,w60,w59,w58,w57,w56,w55,w54,w53,w52,w51,w50,w49,w48,w47,w46,w45,w44,w43,w42,w41,w40,w39,w38,w37,w36,w35,w34,w33,w32,w31,w30,w29,w28,w27,w26,w25,w24,w23,w22,w21,w20,w19,w18,w17,w16,w15,w14,w13,w12,w11,w10,w9,w8,w7,w6,w5,w4,w3}, {w144,w143,w142,w141,w140,w139,w138,w137,w136,w135,w134,w133,w132,w131,w130,w129,w128,w127,w126,w125,w124,w123,w122,w121,w120,w119,w118,w117,w116,w115,w114,w113,w112,w111,w110,w109,w108,w107,w106,w105,w104,w103,w102,w101,w100,w99,w98,w97,w96,w95,w94,w93,w92,w91,w90,w89,w88,w87,w86,w85,w84,w83,w82,w81,w80,w79,w78,w77,w76,w75,w74}, x0_70, {x0_70,x0_69,x0_68,x0_67,x0_66,x0_65,x0_64,x0_63,x0_62,x0_61,x0_60,x0_59,x0_58,x0_57,x0_56,x0_55,x0_54,x0_53,x0_52,x0_51,x0_50,x0_49,x0_48,x0_47,x0_46,x0_45,x0_44,x0_43,x0_42,x0_41,x0_40,x0_39,x0_38,x0_37,x0_36,x0_35,x0_34,x0_33,x0_32,x0_31,x0_30,x0_29,x0_28,x0_27,x0_26,x0_25,x0_24,x0_23,x0_22,x0_21,x0_20,x0_19,x0_18,x0_17,x0_16,x0_15,x0_14,x0_13,x0_12,x0_11,x0_10,x0_9,x0_8,x0_7,x0_6,x0_5,x0_4,x0_3,x0_2,x0_1,x0_0}, {x1_70,x1_69,x1_68,x1_67,x1_66,x1_65,x1_64,x1_63,x1_62,x1_61,x1_60,x1_59,x1_58,x1_57,x1_56,x1_55,x1_54,x1_53,x1_52,x1_51,x1_50,x1_49,x1_48,x1_47,x1_46,x1_45,x1_44,x1_43,x1_42,x1_41,x1_40,x1_39,x1_38,x1_37,x1_36,x1_35,x1_34,x1_33,x1_32,x1_31,x1_30,x1_29,x1_28,x1_27,x1_26,x1_25,x1_24,x1_23,x1_22,x1_21,x1_20,x1_19,x1_18,x1_17,x1_16,x1_15,x1_14,x1_13,x1_12,x1_11,x1_10,x1_9,x1_8,x1_7,x1_6,x1_5,x1_4,x1_3,x1_2,x1_1,x1_0});
    wire w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842;
    sw_m #(.SIZE(71)) sw5({w1771,w1770,w1769,w1768,w1767,w1766,w1765,w1764,w1763,w1762,w1761,w1760,w1759,w1758,w1757,w1756,w1755,w1754,w1753,w1752,w1751,w1750,w1749,w1748,w1747,w1746,w1745,w1744,w1743,w1742,w1741,w1740,w1739,w1738,w1737,w1736,w1735,w1734,w1733,w1732,w1731,w1730,w1729,w1728,w1727,w1726,w1725,w1724,w1723,w1722,w1721,w1720,w1719,w1718,w1717,w1716,w1715,w1714,w1713,w1712,w1711,w1710,w1709,w1708,w1707,w1706,w1705,w1704,w1703,w1702,w1701}, {w1842,w1841,w1840,w1839,w1838,w1837,w1836,w1835,w1834,w1833,w1832,w1831,w1830,w1829,w1828,w1827,w1826,w1825,w1824,w1823,w1822,w1821,w1820,w1819,w1818,w1817,w1816,w1815,w1814,w1813,w1812,w1811,w1810,w1809,w1808,w1807,w1806,w1805,w1804,w1803,w1802,w1801,w1800,w1799,w1798,w1797,w1796,w1795,w1794,w1793,w1792,w1791,w1790,w1789,w1788,w1787,w1786,w1785,w1784,w1783,w1782,w1781,w1780,w1779,w1778,w1777,w1776,w1775,w1774,w1773,w1772}, x12_70, {x12_70,x12_69,x12_68,x12_67,x12_66,x12_65,x12_64,x12_63,x12_62,x12_61,x12_60,x12_59,x12_58,x12_57,x12_56,x12_55,x12_54,x12_53,x12_52,x12_51,x12_50,x12_49,x12_48,x12_47,x12_46,x12_45,x12_44,x12_43,x12_42,x12_41,x12_40,x12_39,x12_38,x12_37,x12_36,x12_35,x12_34,x12_33,x12_32,x12_31,x12_30,x12_29,x12_28,x12_27,x12_26,x12_25,x12_24,x12_23,x12_22,x12_21,x12_20,x12_19,x12_18,x12_17,x12_16,x12_15,x12_14,x12_13,x12_12,x12_11,x12_10,x12_9,x12_8,x12_7,x12_6,x12_5,x12_4,x12_3,x12_2,x12_1,x12_0}, {x13_70,x13_69,x13_68,x13_67,x13_66,x13_65,x13_64,x13_63,x13_62,x13_61,x13_60,x13_59,x13_58,x13_57,x13_56,x13_55,x13_54,x13_53,x13_52,x13_51,x13_50,x13_49,x13_48,x13_47,x13_46,x13_45,x13_44,x13_43,x13_42,x13_41,x13_40,x13_39,x13_38,x13_37,x13_36,x13_35,x13_34,x13_33,x13_32,x13_31,x13_30,x13_29,x13_28,x13_27,x13_26,x13_25,x13_24,x13_23,x13_22,x13_21,x13_20,x13_19,x13_18,x13_17,x13_16,x13_15,x13_14,x13_13,x13_12,x13_11,x13_10,x13_9,x13_8,x13_7,x13_6,x13_5,x13_4,x13_3,x13_2,x13_1,x13_0});
    wire w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710;
    sw_m #(.SIZE(71)) sw6({w639,w638,w637,w636,w635,w634,w633,w632,w631,w630,w629,w628,w627,w626,w625,w624,w623,w622,w621,w620,w619,w618,w617,w616,w615,w614,w613,w612,w611,w610,w609,w608,w607,w606,w605,w604,w603,w602,w601,w600,w599,w598,w597,w596,w595,w594,w593,w592,w591,w590,w589,w588,w587,w586,w585,w584,w583,w582,w581,w580,w579,w578,w577,w576,w575,w574,w573,w572,w571,w570,w569}, {w710,w709,w708,w707,w706,w705,w704,w703,w702,w701,w700,w699,w698,w697,w696,w695,w694,w693,w692,w691,w690,w689,w688,w687,w686,w685,w684,w683,w682,w681,w680,w679,w678,w677,w676,w675,w674,w673,w672,w671,w670,w669,w668,w667,w666,w665,w664,w663,w662,w661,w660,w659,w658,w657,w656,w655,w654,w653,w652,w651,w650,w649,w648,w647,w646,w645,w644,w643,w642,w641,w640}, x4_70, {x4_70,x4_69,x4_68,x4_67,x4_66,x4_65,x4_64,x4_63,x4_62,x4_61,x4_60,x4_59,x4_58,x4_57,x4_56,x4_55,x4_54,x4_53,x4_52,x4_51,x4_50,x4_49,x4_48,x4_47,x4_46,x4_45,x4_44,x4_43,x4_42,x4_41,x4_40,x4_39,x4_38,x4_37,x4_36,x4_35,x4_34,x4_33,x4_32,x4_31,x4_30,x4_29,x4_28,x4_27,x4_26,x4_25,x4_24,x4_23,x4_22,x4_21,x4_20,x4_19,x4_18,x4_17,x4_16,x4_15,x4_14,x4_13,x4_12,x4_11,x4_10,x4_9,x4_8,x4_7,x4_6,x4_5,x4_4,x4_3,x4_2,x4_1,x4_0}, {x5_70,x5_69,x5_68,x5_67,x5_66,x5_65,x5_64,x5_63,x5_62,x5_61,x5_60,x5_59,x5_58,x5_57,x5_56,x5_55,x5_54,x5_53,x5_52,x5_51,x5_50,x5_49,x5_48,x5_47,x5_46,x5_45,x5_44,x5_43,x5_42,x5_41,x5_40,x5_39,x5_38,x5_37,x5_36,x5_35,x5_34,x5_33,x5_32,x5_31,x5_30,x5_29,x5_28,x5_27,x5_26,x5_25,x5_24,x5_23,x5_22,x5_21,x5_20,x5_19,x5_18,x5_17,x5_16,x5_15,x5_14,x5_13,x5_12,x5_11,x5_10,x5_9,x5_8,x5_7,x5_6,x5_5,x5_4,x5_3,x5_2,x5_1,x5_0});
    wire w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276;
    sw_m #(.SIZE(71)) sw7({w1205,w1204,w1203,w1202,w1201,w1200,w1199,w1198,w1197,w1196,w1195,w1194,w1193,w1192,w1191,w1190,w1189,w1188,w1187,w1186,w1185,w1184,w1183,w1182,w1181,w1180,w1179,w1178,w1177,w1176,w1175,w1174,w1173,w1172,w1171,w1170,w1169,w1168,w1167,w1166,w1165,w1164,w1163,w1162,w1161,w1160,w1159,w1158,w1157,w1156,w1155,w1154,w1153,w1152,w1151,w1150,w1149,w1148,w1147,w1146,w1145,w1144,w1143,w1142,w1141,w1140,w1139,w1138,w1137,w1136,w1135}, {w1276,w1275,w1274,w1273,w1272,w1271,w1270,w1269,w1268,w1267,w1266,w1265,w1264,w1263,w1262,w1261,w1260,w1259,w1258,w1257,w1256,w1255,w1254,w1253,w1252,w1251,w1250,w1249,w1248,w1247,w1246,w1245,w1244,w1243,w1242,w1241,w1240,w1239,w1238,w1237,w1236,w1235,w1234,w1233,w1232,w1231,w1230,w1229,w1228,w1227,w1226,w1225,w1224,w1223,w1222,w1221,w1220,w1219,w1218,w1217,w1216,w1215,w1214,w1213,w1212,w1211,w1210,w1209,w1208,w1207,w1206}, x8_70, {x8_70,x8_69,x8_68,x8_67,x8_66,x8_65,x8_64,x8_63,x8_62,x8_61,x8_60,x8_59,x8_58,x8_57,x8_56,x8_55,x8_54,x8_53,x8_52,x8_51,x8_50,x8_49,x8_48,x8_47,x8_46,x8_45,x8_44,x8_43,x8_42,x8_41,x8_40,x8_39,x8_38,x8_37,x8_36,x8_35,x8_34,x8_33,x8_32,x8_31,x8_30,x8_29,x8_28,x8_27,x8_26,x8_25,x8_24,x8_23,x8_22,x8_21,x8_20,x8_19,x8_18,x8_17,x8_16,x8_15,x8_14,x8_13,x8_12,x8_11,x8_10,x8_9,x8_8,x8_7,x8_6,x8_5,x8_4,x8_3,x8_2,x8_1,x8_0}, {x9_70,x9_69,x9_68,x9_67,x9_66,x9_65,x9_64,x9_63,x9_62,x9_61,x9_60,x9_59,x9_58,x9_57,x9_56,x9_55,x9_54,x9_53,x9_52,x9_51,x9_50,x9_49,x9_48,x9_47,x9_46,x9_45,x9_44,x9_43,x9_42,x9_41,x9_40,x9_39,x9_38,x9_37,x9_36,x9_35,x9_34,x9_33,x9_32,x9_31,x9_30,x9_29,x9_28,x9_27,x9_26,x9_25,x9_24,x9_23,x9_22,x9_21,x9_20,x9_19,x9_18,x9_17,x9_16,x9_15,x9_14,x9_13,x9_12,x9_11,x9_10,x9_9,x9_8,x9_7,x9_6,x9_5,x9_4,x9_3,x9_2,x9_1,x9_0});
    wire w2;
    xor xor8(w2, x0_70, w1);
    wire w1700;
    xor xor9(w1700, x12_70, w1699);
    wire w568;
    xor xor10(w568, x4_70, w567);
    wire w1134;
    xor xor11(w1134, x8_70, w1133);
    wire w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418;
    sw_m #(.SIZE(71)) sw12({w1347,w1346,w1345,w1344,w1343,w1342,w1341,w1340,w1339,w1338,w1337,w1336,w1335,w1334,w1333,w1332,w1331,w1330,w1329,w1328,w1327,w1326,w1325,w1324,w1323,w1322,w1321,w1320,w1319,w1318,w1317,w1316,w1315,w1314,w1313,w1312,w1311,w1310,w1309,w1308,w1307,w1306,w1305,w1304,w1303,w1302,w1301,w1300,w1299,w1298,w1297,w1296,w1295,w1294,w1293,w1292,w1291,w1290,w1289,w1288,w1287,w1286,w1285,w1284,w1283,w1282,w1281,w1280,w1279,w1278,w1277}, {w1418,w1417,w1416,w1415,w1414,w1413,w1412,w1411,w1410,w1409,w1408,w1407,w1406,w1405,w1404,w1403,w1402,w1401,w1400,w1399,w1398,w1397,w1396,w1395,w1394,w1393,w1392,w1391,w1390,w1389,w1388,w1387,w1386,w1385,w1384,w1383,w1382,w1381,w1380,w1379,w1378,w1377,w1376,w1375,w1374,w1373,w1372,w1371,w1370,w1369,w1368,w1367,w1366,w1365,w1364,w1363,w1362,w1361,w1360,w1359,w1358,w1357,w1356,w1355,w1354,w1353,w1352,w1351,w1350,w1349,w1348}, w1134, {x10_70,x10_69,x10_68,x10_67,x10_66,x10_65,x10_64,x10_63,x10_62,x10_61,x10_60,x10_59,x10_58,x10_57,x10_56,x10_55,x10_54,x10_53,x10_52,x10_51,x10_50,x10_49,x10_48,x10_47,x10_46,x10_45,x10_44,x10_43,x10_42,x10_41,x10_40,x10_39,x10_38,x10_37,x10_36,x10_35,x10_34,x10_33,x10_32,x10_31,x10_30,x10_29,x10_28,x10_27,x10_26,x10_25,x10_24,x10_23,x10_22,x10_21,x10_20,x10_19,x10_18,x10_17,x10_16,x10_15,x10_14,x10_13,x10_12,x10_11,x10_10,x10_9,x10_8,x10_7,x10_6,x10_5,x10_4,x10_3,x10_2,x10_1,x10_0}, {x11_70,x11_69,x11_68,x11_67,x11_66,x11_65,x11_64,x11_63,x11_62,x11_61,x11_60,x11_59,x11_58,x11_57,x11_56,x11_55,x11_54,x11_53,x11_52,x11_51,x11_50,x11_49,x11_48,x11_47,x11_46,x11_45,x11_44,x11_43,x11_42,x11_41,x11_40,x11_39,x11_38,x11_37,x11_36,x11_35,x11_34,x11_33,x11_32,x11_31,x11_30,x11_29,x11_28,x11_27,x11_26,x11_25,x11_24,x11_23,x11_22,x11_21,x11_20,x11_19,x11_18,x11_17,x11_16,x11_15,x11_14,x11_13,x11_12,x11_11,x11_10,x11_9,x11_8,x11_7,x11_6,x11_5,x11_4,x11_3,x11_2,x11_1,x11_0});
    wire w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984;
    sw_m #(.SIZE(71)) sw13({w1913,w1912,w1911,w1910,w1909,w1908,w1907,w1906,w1905,w1904,w1903,w1902,w1901,w1900,w1899,w1898,w1897,w1896,w1895,w1894,w1893,w1892,w1891,w1890,w1889,w1888,w1887,w1886,w1885,w1884,w1883,w1882,w1881,w1880,w1879,w1878,w1877,w1876,w1875,w1874,w1873,w1872,w1871,w1870,w1869,w1868,w1867,w1866,w1865,w1864,w1863,w1862,w1861,w1860,w1859,w1858,w1857,w1856,w1855,w1854,w1853,w1852,w1851,w1850,w1849,w1848,w1847,w1846,w1845,w1844,w1843}, {w1984,w1983,w1982,w1981,w1980,w1979,w1978,w1977,w1976,w1975,w1974,w1973,w1972,w1971,w1970,w1969,w1968,w1967,w1966,w1965,w1964,w1963,w1962,w1961,w1960,w1959,w1958,w1957,w1956,w1955,w1954,w1953,w1952,w1951,w1950,w1949,w1948,w1947,w1946,w1945,w1944,w1943,w1942,w1941,w1940,w1939,w1938,w1937,w1936,w1935,w1934,w1933,w1932,w1931,w1930,w1929,w1928,w1927,w1926,w1925,w1924,w1923,w1922,w1921,w1920,w1919,w1918,w1917,w1916,w1915,w1914}, w1700, {x14_70,x14_69,x14_68,x14_67,x14_66,x14_65,x14_64,x14_63,x14_62,x14_61,x14_60,x14_59,x14_58,x14_57,x14_56,x14_55,x14_54,x14_53,x14_52,x14_51,x14_50,x14_49,x14_48,x14_47,x14_46,x14_45,x14_44,x14_43,x14_42,x14_41,x14_40,x14_39,x14_38,x14_37,x14_36,x14_35,x14_34,x14_33,x14_32,x14_31,x14_30,x14_29,x14_28,x14_27,x14_26,x14_25,x14_24,x14_23,x14_22,x14_21,x14_20,x14_19,x14_18,x14_17,x14_16,x14_15,x14_14,x14_13,x14_12,x14_11,x14_10,x14_9,x14_8,x14_7,x14_6,x14_5,x14_4,x14_3,x14_2,x14_1,x14_0}, {x15_70,x15_69,x15_68,x15_67,x15_66,x15_65,x15_64,x15_63,x15_62,x15_61,x15_60,x15_59,x15_58,x15_57,x15_56,x15_55,x15_54,x15_53,x15_52,x15_51,x15_50,x15_49,x15_48,x15_47,x15_46,x15_45,x15_44,x15_43,x15_42,x15_41,x15_40,x15_39,x15_38,x15_37,x15_36,x15_35,x15_34,x15_33,x15_32,x15_31,x15_30,x15_29,x15_28,x15_27,x15_26,x15_25,x15_24,x15_23,x15_22,x15_21,x15_20,x15_19,x15_18,x15_17,x15_16,x15_15,x15_14,x15_13,x15_12,x15_11,x15_10,x15_9,x15_8,x15_7,x15_6,x15_5,x15_4,x15_3,x15_2,x15_1,x15_0});
    wire w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286;
    sw_m #(.SIZE(71)) sw14({w215,w214,w213,w212,w211,w210,w209,w208,w207,w206,w205,w204,w203,w202,w201,w200,w199,w198,w197,w196,w195,w194,w193,w192,w191,w190,w189,w188,w187,w186,w185,w184,w183,w182,w181,w180,w179,w178,w177,w176,w175,w174,w173,w172,w171,w170,w169,w168,w167,w166,w165,w164,w163,w162,w161,w160,w159,w158,w157,w156,w155,w154,w153,w152,w151,w150,w149,w148,w147,w146,w145}, {w286,w285,w284,w283,w282,w281,w280,w279,w278,w277,w276,w275,w274,w273,w272,w271,w270,w269,w268,w267,w266,w265,w264,w263,w262,w261,w260,w259,w258,w257,w256,w255,w254,w253,w252,w251,w250,w249,w248,w247,w246,w245,w244,w243,w242,w241,w240,w239,w238,w237,w236,w235,w234,w233,w232,w231,w230,w229,w228,w227,w226,w225,w224,w223,w222,w221,w220,w219,w218,w217,w216}, w2, {x2_70,x2_69,x2_68,x2_67,x2_66,x2_65,x2_64,x2_63,x2_62,x2_61,x2_60,x2_59,x2_58,x2_57,x2_56,x2_55,x2_54,x2_53,x2_52,x2_51,x2_50,x2_49,x2_48,x2_47,x2_46,x2_45,x2_44,x2_43,x2_42,x2_41,x2_40,x2_39,x2_38,x2_37,x2_36,x2_35,x2_34,x2_33,x2_32,x2_31,x2_30,x2_29,x2_28,x2_27,x2_26,x2_25,x2_24,x2_23,x2_22,x2_21,x2_20,x2_19,x2_18,x2_17,x2_16,x2_15,x2_14,x2_13,x2_12,x2_11,x2_10,x2_9,x2_8,x2_7,x2_6,x2_5,x2_4,x2_3,x2_2,x2_1,x2_0}, {x3_70,x3_69,x3_68,x3_67,x3_66,x3_65,x3_64,x3_63,x3_62,x3_61,x3_60,x3_59,x3_58,x3_57,x3_56,x3_55,x3_54,x3_53,x3_52,x3_51,x3_50,x3_49,x3_48,x3_47,x3_46,x3_45,x3_44,x3_43,x3_42,x3_41,x3_40,x3_39,x3_38,x3_37,x3_36,x3_35,x3_34,x3_33,x3_32,x3_31,x3_30,x3_29,x3_28,x3_27,x3_26,x3_25,x3_24,x3_23,x3_22,x3_21,x3_20,x3_19,x3_18,x3_17,x3_16,x3_15,x3_14,x3_13,x3_12,x3_11,x3_10,x3_9,x3_8,x3_7,x3_6,x3_5,x3_4,x3_3,x3_2,x3_1,x3_0});
    wire w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852;
    sw_m #(.SIZE(71)) sw15({w781,w780,w779,w778,w777,w776,w775,w774,w773,w772,w771,w770,w769,w768,w767,w766,w765,w764,w763,w762,w761,w760,w759,w758,w757,w756,w755,w754,w753,w752,w751,w750,w749,w748,w747,w746,w745,w744,w743,w742,w741,w740,w739,w738,w737,w736,w735,w734,w733,w732,w731,w730,w729,w728,w727,w726,w725,w724,w723,w722,w721,w720,w719,w718,w717,w716,w715,w714,w713,w712,w711}, {w852,w851,w850,w849,w848,w847,w846,w845,w844,w843,w842,w841,w840,w839,w838,w837,w836,w835,w834,w833,w832,w831,w830,w829,w828,w827,w826,w825,w824,w823,w822,w821,w820,w819,w818,w817,w816,w815,w814,w813,w812,w811,w810,w809,w808,w807,w806,w805,w804,w803,w802,w801,w800,w799,w798,w797,w796,w795,w794,w793,w792,w791,w790,w789,w788,w787,w786,w785,w784,w783,w782}, w568, {x6_70,x6_69,x6_68,x6_67,x6_66,x6_65,x6_64,x6_63,x6_62,x6_61,x6_60,x6_59,x6_58,x6_57,x6_56,x6_55,x6_54,x6_53,x6_52,x6_51,x6_50,x6_49,x6_48,x6_47,x6_46,x6_45,x6_44,x6_43,x6_42,x6_41,x6_40,x6_39,x6_38,x6_37,x6_36,x6_35,x6_34,x6_33,x6_32,x6_31,x6_30,x6_29,x6_28,x6_27,x6_26,x6_25,x6_24,x6_23,x6_22,x6_21,x6_20,x6_19,x6_18,x6_17,x6_16,x6_15,x6_14,x6_13,x6_12,x6_11,x6_10,x6_9,x6_8,x6_7,x6_6,x6_5,x6_4,x6_3,x6_2,x6_1,x6_0}, {x7_70,x7_69,x7_68,x7_67,x7_66,x7_65,x7_64,x7_63,x7_62,x7_61,x7_60,x7_59,x7_58,x7_57,x7_56,x7_55,x7_54,x7_53,x7_52,x7_51,x7_50,x7_49,x7_48,x7_47,x7_46,x7_45,x7_44,x7_43,x7_42,x7_41,x7_40,x7_39,x7_38,x7_37,x7_36,x7_35,x7_34,x7_33,x7_32,x7_31,x7_30,x7_29,x7_28,x7_27,x7_26,x7_25,x7_24,x7_23,x7_22,x7_21,x7_20,x7_19,x7_18,x7_17,x7_16,x7_15,x7_14,x7_13,x7_12,x7_11,x7_10,x7_9,x7_8,x7_7,x7_6,x7_5,x7_4,x7_3,x7_2,x7_1,x7_0});
    sw_m #(.SIZE(70)) sw16({w1488,w1487,w1486,w1485,w1484,w1483,w1482,w1481,w1480,w1479,w1478,w1477,w1476,w1475,w1474,w1473,w1472,w1471,w1470,w1469,w1468,w1467,w1466,w1465,w1464,w1463,w1462,w1461,w1460,w1459,w1458,w1457,w1456,w1455,w1454,w1453,w1452,w1451,w1450,w1449,w1448,w1447,w1446,w1445,w1444,w1443,w1442,w1441,w1440,w1439,w1438,w1437,w1436,w1435,w1434,w1433,w1432,w1431,w1430,w1429,w1428,w1427,w1426,w1425,w1424,w1423,w1422,w1421,w1420,w1419}, {w1558,w1557,w1556,w1555,w1554,w1553,w1552,w1551,w1550,w1549,w1548,w1547,w1546,w1545,w1544,w1543,w1542,w1541,w1540,w1539,w1538,w1537,w1536,w1535,w1534,w1533,w1532,w1531,w1530,w1529,w1528,w1527,w1526,w1525,w1524,w1523,w1522,w1521,w1520,w1519,w1518,w1517,w1516,w1515,w1514,w1513,w1512,w1511,w1510,w1509,w1508,w1507,w1506,w1505,w1504,w1503,w1502,w1501,w1500,w1499,w1498,w1497,w1496,w1495,w1494,w1493,w1492,w1491,w1490,w1489}, w1205, {w1204,w1203,w1202,w1201,w1200,w1199,w1198,w1197,w1196,w1195,w1194,w1193,w1192,w1191,w1190,w1189,w1188,w1187,w1186,w1185,w1184,w1183,w1182,w1181,w1180,w1179,w1178,w1177,w1176,w1175,w1174,w1173,w1172,w1171,w1170,w1169,w1168,w1167,w1166,w1165,w1164,w1163,w1162,w1161,w1160,w1159,w1158,w1157,w1156,w1155,w1154,w1153,w1152,w1151,w1150,w1149,w1148,w1147,w1146,w1145,w1144,w1143,w1142,w1141,w1140,w1139,w1138,w1137,w1136,w1135}, {w1346,w1345,w1344,w1343,w1342,w1341,w1340,w1339,w1338,w1337,w1336,w1335,w1334,w1333,w1332,w1331,w1330,w1329,w1328,w1327,w1326,w1325,w1324,w1323,w1322,w1321,w1320,w1319,w1318,w1317,w1316,w1315,w1314,w1313,w1312,w1311,w1310,w1309,w1308,w1307,w1306,w1305,w1304,w1303,w1302,w1301,w1300,w1299,w1298,w1297,w1296,w1295,w1294,w1293,w1292,w1291,w1290,w1289,w1288,w1287,w1286,w1285,w1284,w1283,w1282,w1281,w1280,w1279,w1278,w1277});
    sw_m #(.SIZE(70)) sw17({w1628,w1627,w1626,w1625,w1624,w1623,w1622,w1621,w1620,w1619,w1618,w1617,w1616,w1615,w1614,w1613,w1612,w1611,w1610,w1609,w1608,w1607,w1606,w1605,w1604,w1603,w1602,w1601,w1600,w1599,w1598,w1597,w1596,w1595,w1594,w1593,w1592,w1591,w1590,w1589,w1588,w1587,w1586,w1585,w1584,w1583,w1582,w1581,w1580,w1579,w1578,w1577,w1576,w1575,w1574,w1573,w1572,w1571,w1570,w1569,w1568,w1567,w1566,w1565,w1564,w1563,w1562,w1561,w1560,w1559}, {w1698,w1697,w1696,w1695,w1694,w1693,w1692,w1691,w1690,w1689,w1688,w1687,w1686,w1685,w1684,w1683,w1682,w1681,w1680,w1679,w1678,w1677,w1676,w1675,w1674,w1673,w1672,w1671,w1670,w1669,w1668,w1667,w1666,w1665,w1664,w1663,w1662,w1661,w1660,w1659,w1658,w1657,w1656,w1655,w1654,w1653,w1652,w1651,w1650,w1649,w1648,w1647,w1646,w1645,w1644,w1643,w1642,w1641,w1640,w1639,w1638,w1637,w1636,w1635,w1634,w1633,w1632,w1631,w1630,w1629}, w1276, {w1275,w1274,w1273,w1272,w1271,w1270,w1269,w1268,w1267,w1266,w1265,w1264,w1263,w1262,w1261,w1260,w1259,w1258,w1257,w1256,w1255,w1254,w1253,w1252,w1251,w1250,w1249,w1248,w1247,w1246,w1245,w1244,w1243,w1242,w1241,w1240,w1239,w1238,w1237,w1236,w1235,w1234,w1233,w1232,w1231,w1230,w1229,w1228,w1227,w1226,w1225,w1224,w1223,w1222,w1221,w1220,w1219,w1218,w1217,w1216,w1215,w1214,w1213,w1212,w1211,w1210,w1209,w1208,w1207,w1206}, {w1417,w1416,w1415,w1414,w1413,w1412,w1411,w1410,w1409,w1408,w1407,w1406,w1405,w1404,w1403,w1402,w1401,w1400,w1399,w1398,w1397,w1396,w1395,w1394,w1393,w1392,w1391,w1390,w1389,w1388,w1387,w1386,w1385,w1384,w1383,w1382,w1381,w1380,w1379,w1378,w1377,w1376,w1375,w1374,w1373,w1372,w1371,w1370,w1369,w1368,w1367,w1366,w1365,w1364,w1363,w1362,w1361,w1360,w1359,w1358,w1357,w1356,w1355,w1354,w1353,w1352,w1351,w1350,w1349,w1348});
    sw_m #(.SIZE(70)) sw18({w496,w495,w494,w493,w492,w491,w490,w489,w488,w487,w486,w485,w484,w483,w482,w481,w480,w479,w478,w477,w476,w475,w474,w473,w472,w471,w470,w469,w468,w467,w466,w465,w464,w463,w462,w461,w460,w459,w458,w457,w456,w455,w454,w453,w452,w451,w450,w449,w448,w447,w446,w445,w444,w443,w442,w441,w440,w439,w438,w437,w436,w435,w434,w433,w432,w431,w430,w429,w428,w427}, {w566,w565,w564,w563,w562,w561,w560,w559,w558,w557,w556,w555,w554,w553,w552,w551,w550,w549,w548,w547,w546,w545,w544,w543,w542,w541,w540,w539,w538,w537,w536,w535,w534,w533,w532,w531,w530,w529,w528,w527,w526,w525,w524,w523,w522,w521,w520,w519,w518,w517,w516,w515,w514,w513,w512,w511,w510,w509,w508,w507,w506,w505,w504,w503,w502,w501,w500,w499,w498,w497}, w144, {w143,w142,w141,w140,w139,w138,w137,w136,w135,w134,w133,w132,w131,w130,w129,w128,w127,w126,w125,w124,w123,w122,w121,w120,w119,w118,w117,w116,w115,w114,w113,w112,w111,w110,w109,w108,w107,w106,w105,w104,w103,w102,w101,w100,w99,w98,w97,w96,w95,w94,w93,w92,w91,w90,w89,w88,w87,w86,w85,w84,w83,w82,w81,w80,w79,w78,w77,w76,w75,w74}, {w285,w284,w283,w282,w281,w280,w279,w278,w277,w276,w275,w274,w273,w272,w271,w270,w269,w268,w267,w266,w265,w264,w263,w262,w261,w260,w259,w258,w257,w256,w255,w254,w253,w252,w251,w250,w249,w248,w247,w246,w245,w244,w243,w242,w241,w240,w239,w238,w237,w236,w235,w234,w233,w232,w231,w230,w229,w228,w227,w226,w225,w224,w223,w222,w221,w220,w219,w218,w217,w216});
    sw_m #(.SIZE(70)) sw19({w2054,w2053,w2052,w2051,w2050,w2049,w2048,w2047,w2046,w2045,w2044,w2043,w2042,w2041,w2040,w2039,w2038,w2037,w2036,w2035,w2034,w2033,w2032,w2031,w2030,w2029,w2028,w2027,w2026,w2025,w2024,w2023,w2022,w2021,w2020,w2019,w2018,w2017,w2016,w2015,w2014,w2013,w2012,w2011,w2010,w2009,w2008,w2007,w2006,w2005,w2004,w2003,w2002,w2001,w2000,w1999,w1998,w1997,w1996,w1995,w1994,w1993,w1992,w1991,w1990,w1989,w1988,w1987,w1986,w1985}, {w2124,w2123,w2122,w2121,w2120,w2119,w2118,w2117,w2116,w2115,w2114,w2113,w2112,w2111,w2110,w2109,w2108,w2107,w2106,w2105,w2104,w2103,w2102,w2101,w2100,w2099,w2098,w2097,w2096,w2095,w2094,w2093,w2092,w2091,w2090,w2089,w2088,w2087,w2086,w2085,w2084,w2083,w2082,w2081,w2080,w2079,w2078,w2077,w2076,w2075,w2074,w2073,w2072,w2071,w2070,w2069,w2068,w2067,w2066,w2065,w2064,w2063,w2062,w2061,w2060,w2059,w2058,w2057,w2056,w2055}, w1771, {w1770,w1769,w1768,w1767,w1766,w1765,w1764,w1763,w1762,w1761,w1760,w1759,w1758,w1757,w1756,w1755,w1754,w1753,w1752,w1751,w1750,w1749,w1748,w1747,w1746,w1745,w1744,w1743,w1742,w1741,w1740,w1739,w1738,w1737,w1736,w1735,w1734,w1733,w1732,w1731,w1730,w1729,w1728,w1727,w1726,w1725,w1724,w1723,w1722,w1721,w1720,w1719,w1718,w1717,w1716,w1715,w1714,w1713,w1712,w1711,w1710,w1709,w1708,w1707,w1706,w1705,w1704,w1703,w1702,w1701}, {w1912,w1911,w1910,w1909,w1908,w1907,w1906,w1905,w1904,w1903,w1902,w1901,w1900,w1899,w1898,w1897,w1896,w1895,w1894,w1893,w1892,w1891,w1890,w1889,w1888,w1887,w1886,w1885,w1884,w1883,w1882,w1881,w1880,w1879,w1878,w1877,w1876,w1875,w1874,w1873,w1872,w1871,w1870,w1869,w1868,w1867,w1866,w1865,w1864,w1863,w1862,w1861,w1860,w1859,w1858,w1857,w1856,w1855,w1854,w1853,w1852,w1851,w1850,w1849,w1848,w1847,w1846,w1845,w1844,w1843});
    sw_m #(.SIZE(70)) sw20({w2194,w2193,w2192,w2191,w2190,w2189,w2188,w2187,w2186,w2185,w2184,w2183,w2182,w2181,w2180,w2179,w2178,w2177,w2176,w2175,w2174,w2173,w2172,w2171,w2170,w2169,w2168,w2167,w2166,w2165,w2164,w2163,w2162,w2161,w2160,w2159,w2158,w2157,w2156,w2155,w2154,w2153,w2152,w2151,w2150,w2149,w2148,w2147,w2146,w2145,w2144,w2143,w2142,w2141,w2140,w2139,w2138,w2137,w2136,w2135,w2134,w2133,w2132,w2131,w2130,w2129,w2128,w2127,w2126,w2125}, {w2264,w2263,w2262,w2261,w2260,w2259,w2258,w2257,w2256,w2255,w2254,w2253,w2252,w2251,w2250,w2249,w2248,w2247,w2246,w2245,w2244,w2243,w2242,w2241,w2240,w2239,w2238,w2237,w2236,w2235,w2234,w2233,w2232,w2231,w2230,w2229,w2228,w2227,w2226,w2225,w2224,w2223,w2222,w2221,w2220,w2219,w2218,w2217,w2216,w2215,w2214,w2213,w2212,w2211,w2210,w2209,w2208,w2207,w2206,w2205,w2204,w2203,w2202,w2201,w2200,w2199,w2198,w2197,w2196,w2195}, w1842, {w1841,w1840,w1839,w1838,w1837,w1836,w1835,w1834,w1833,w1832,w1831,w1830,w1829,w1828,w1827,w1826,w1825,w1824,w1823,w1822,w1821,w1820,w1819,w1818,w1817,w1816,w1815,w1814,w1813,w1812,w1811,w1810,w1809,w1808,w1807,w1806,w1805,w1804,w1803,w1802,w1801,w1800,w1799,w1798,w1797,w1796,w1795,w1794,w1793,w1792,w1791,w1790,w1789,w1788,w1787,w1786,w1785,w1784,w1783,w1782,w1781,w1780,w1779,w1778,w1777,w1776,w1775,w1774,w1773,w1772}, {w1983,w1982,w1981,w1980,w1979,w1978,w1977,w1976,w1975,w1974,w1973,w1972,w1971,w1970,w1969,w1968,w1967,w1966,w1965,w1964,w1963,w1962,w1961,w1960,w1959,w1958,w1957,w1956,w1955,w1954,w1953,w1952,w1951,w1950,w1949,w1948,w1947,w1946,w1945,w1944,w1943,w1942,w1941,w1940,w1939,w1938,w1937,w1936,w1935,w1934,w1933,w1932,w1931,w1930,w1929,w1928,w1927,w1926,w1925,w1924,w1923,w1922,w1921,w1920,w1919,w1918,w1917,w1916,w1915,w1914});
    sw_m #(.SIZE(70)) sw21({w922,w921,w920,w919,w918,w917,w916,w915,w914,w913,w912,w911,w910,w909,w908,w907,w906,w905,w904,w903,w902,w901,w900,w899,w898,w897,w896,w895,w894,w893,w892,w891,w890,w889,w888,w887,w886,w885,w884,w883,w882,w881,w880,w879,w878,w877,w876,w875,w874,w873,w872,w871,w870,w869,w868,w867,w866,w865,w864,w863,w862,w861,w860,w859,w858,w857,w856,w855,w854,w853}, {w992,w991,w990,w989,w988,w987,w986,w985,w984,w983,w982,w981,w980,w979,w978,w977,w976,w975,w974,w973,w972,w971,w970,w969,w968,w967,w966,w965,w964,w963,w962,w961,w960,w959,w958,w957,w956,w955,w954,w953,w952,w951,w950,w949,w948,w947,w946,w945,w944,w943,w942,w941,w940,w939,w938,w937,w936,w935,w934,w933,w932,w931,w930,w929,w928,w927,w926,w925,w924,w923}, w639, {w638,w637,w636,w635,w634,w633,w632,w631,w630,w629,w628,w627,w626,w625,w624,w623,w622,w621,w620,w619,w618,w617,w616,w615,w614,w613,w612,w611,w610,w609,w608,w607,w606,w605,w604,w603,w602,w601,w600,w599,w598,w597,w596,w595,w594,w593,w592,w591,w590,w589,w588,w587,w586,w585,w584,w583,w582,w581,w580,w579,w578,w577,w576,w575,w574,w573,w572,w571,w570,w569}, {w780,w779,w778,w777,w776,w775,w774,w773,w772,w771,w770,w769,w768,w767,w766,w765,w764,w763,w762,w761,w760,w759,w758,w757,w756,w755,w754,w753,w752,w751,w750,w749,w748,w747,w746,w745,w744,w743,w742,w741,w740,w739,w738,w737,w736,w735,w734,w733,w732,w731,w730,w729,w728,w727,w726,w725,w724,w723,w722,w721,w720,w719,w718,w717,w716,w715,w714,w713,w712,w711});
    sw_m #(.SIZE(70)) sw22({w1062,w1061,w1060,w1059,w1058,w1057,w1056,w1055,w1054,w1053,w1052,w1051,w1050,w1049,w1048,w1047,w1046,w1045,w1044,w1043,w1042,w1041,w1040,w1039,w1038,w1037,w1036,w1035,w1034,w1033,w1032,w1031,w1030,w1029,w1028,w1027,w1026,w1025,w1024,w1023,w1022,w1021,w1020,w1019,w1018,w1017,w1016,w1015,w1014,w1013,w1012,w1011,w1010,w1009,w1008,w1007,w1006,w1005,w1004,w1003,w1002,w1001,w1000,w999,w998,w997,w996,w995,w994,w993}, {w1132,w1131,w1130,w1129,w1128,w1127,w1126,w1125,w1124,w1123,w1122,w1121,w1120,w1119,w1118,w1117,w1116,w1115,w1114,w1113,w1112,w1111,w1110,w1109,w1108,w1107,w1106,w1105,w1104,w1103,w1102,w1101,w1100,w1099,w1098,w1097,w1096,w1095,w1094,w1093,w1092,w1091,w1090,w1089,w1088,w1087,w1086,w1085,w1084,w1083,w1082,w1081,w1080,w1079,w1078,w1077,w1076,w1075,w1074,w1073,w1072,w1071,w1070,w1069,w1068,w1067,w1066,w1065,w1064,w1063}, w710, {w709,w708,w707,w706,w705,w704,w703,w702,w701,w700,w699,w698,w697,w696,w695,w694,w693,w692,w691,w690,w689,w688,w687,w686,w685,w684,w683,w682,w681,w680,w679,w678,w677,w676,w675,w674,w673,w672,w671,w670,w669,w668,w667,w666,w665,w664,w663,w662,w661,w660,w659,w658,w657,w656,w655,w654,w653,w652,w651,w650,w649,w648,w647,w646,w645,w644,w643,w642,w641,w640}, {w851,w850,w849,w848,w847,w846,w845,w844,w843,w842,w841,w840,w839,w838,w837,w836,w835,w834,w833,w832,w831,w830,w829,w828,w827,w826,w825,w824,w823,w822,w821,w820,w819,w818,w817,w816,w815,w814,w813,w812,w811,w810,w809,w808,w807,w806,w805,w804,w803,w802,w801,w800,w799,w798,w797,w796,w795,w794,w793,w792,w791,w790,w789,w788,w787,w786,w785,w784,w783,w782});
    sw_m #(.SIZE(70)) sw23({w356,w355,w354,w353,w352,w351,w350,w349,w348,w347,w346,w345,w344,w343,w342,w341,w340,w339,w338,w337,w336,w335,w334,w333,w332,w331,w330,w329,w328,w327,w326,w325,w324,w323,w322,w321,w320,w319,w318,w317,w316,w315,w314,w313,w312,w311,w310,w309,w308,w307,w306,w305,w304,w303,w302,w301,w300,w299,w298,w297,w296,w295,w294,w293,w292,w291,w290,w289,w288,w287}, {w426,w425,w424,w423,w422,w421,w420,w419,w418,w417,w416,w415,w414,w413,w412,w411,w410,w409,w408,w407,w406,w405,w404,w403,w402,w401,w400,w399,w398,w397,w396,w395,w394,w393,w392,w391,w390,w389,w388,w387,w386,w385,w384,w383,w382,w381,w380,w379,w378,w377,w376,w375,w374,w373,w372,w371,w370,w369,w368,w367,w366,w365,w364,w363,w362,w361,w360,w359,w358,w357}, w73, {w72,w71,w70,w69,w68,w67,w66,w65,w64,w63,w62,w61,w60,w59,w58,w57,w56,w55,w54,w53,w52,w51,w50,w49,w48,w47,w46,w45,w44,w43,w42,w41,w40,w39,w38,w37,w36,w35,w34,w33,w32,w31,w30,w29,w28,w27,w26,w25,w24,w23,w22,w21,w20,w19,w18,w17,w16,w15,w14,w13,w12,w11,w10,w9,w8,w7,w6,w5,w4,w3}, {w214,w213,w212,w211,w210,w209,w208,w207,w206,w205,w204,w203,w202,w201,w200,w199,w198,w197,w196,w195,w194,w193,w192,w191,w190,w189,w188,w187,w186,w185,w184,w183,w182,w181,w180,w179,w178,w177,w176,w175,w174,w173,w172,w171,w170,w169,w168,w167,w166,w165,w164,w163,w162,w161,w160,w159,w158,w157,w156,w155,w154,w153,w152,w151,w150,w149,w148,w147,w146,w145});
endmodule
