`default_nettype none

module TNT_BIN_HC0_JaSJ17_68_16_0_pipelined(input wire clock, message_interface_nonblocking.producer out0, message_interface_nonblocking.producer out1, message_interface_nonblocking.producer out2, message_interface_nonblocking.producer out3, message_interface_nonblocking.producer out4, message_interface_nonblocking.producer out5, message_interface_nonblocking.producer out6, message_interface_nonblocking.producer out7, message_interface_nonblocking.producer out8, message_interface_nonblocking.producer out9, message_interface_nonblocking.producer out10, message_interface_nonblocking.producer out11, message_interface_nonblocking.producer out12, message_interface_nonblocking.producer out13, message_interface_nonblocking.producer out14, message_interface_nonblocking.producer out15, message_interface_nonblocking.consumer in0, message_interface_nonblocking.consumer in1, message_interface_nonblocking.consumer in2, message_interface_nonblocking.consumer in3, message_interface_nonblocking.consumer in4, message_interface_nonblocking.consumer in5, message_interface_nonblocking.consumer in6, message_interface_nonblocking.consumer in7, message_interface_nonblocking.consumer in8, message_interface_nonblocking.consumer in9, message_interface_nonblocking.consumer in10, message_interface_nonblocking.consumer in11, message_interface_nonblocking.consumer in12, message_interface_nonblocking.consumer in13, message_interface_nonblocking.consumer in14, message_interface_nonblocking.consumer in15);
wire [72:0] internal_in0;
wire [72:0] internal_in1;
wire [72:0] internal_in2;
wire [72:0] internal_in3;
wire [72:0] internal_in4;
wire [72:0] internal_in5;
wire [72:0] internal_in6;
wire [72:0] internal_in7;
wire [72:0] internal_in8;
wire [72:0] internal_in9;
wire [72:0] internal_in10;
wire [72:0] internal_in11;
wire [72:0] internal_in12;
wire [72:0] internal_in13;
wire [72:0] internal_in14;
wire [72:0] internal_in15;
wire [69:0] internal_out0;
wire [69:0] internal_out1;
wire [69:0] internal_out2;
wire [69:0] internal_out3;
wire [69:0] internal_out4;
wire [69:0] internal_out5;
wire [69:0] internal_out6;
wire [69:0] internal_out7;
wire [69:0] internal_out8;
wire [69:0] internal_out9;
wire [69:0] internal_out10;
wire [69:0] internal_out11;
wire [69:0] internal_out12;
wire [69:0] internal_out13;
wire [69:0] internal_out14;
wire [69:0] internal_out15;
wire [72:0] between_0_0;
wire [72:0] between_1_0;
wire [72:0] between_2_0;
wire [72:0] between_3_0;
wire [72:0] between_4_0;
wire [72:0] between_5_0;
wire [72:0] between_6_0;
wire [72:0] between_7_0;
wire [72:0] between_8_0;
wire [72:0] between_9_0;
wire [72:0] between_10_0;
wire [72:0] between_11_0;
wire [72:0] between_12_0;
wire [72:0] between_13_0;
wire [72:0] between_14_0;
wire [72:0] between_15_0;
wire [72:0] between_0_1;
wire [72:0] between_1_1;
wire [72:0] between_2_1;
wire [72:0] between_3_1;
wire [72:0] between_4_1;
wire [72:0] between_5_1;
wire [72:0] between_6_1;
wire [72:0] between_7_1;
wire [72:0] between_8_1;
wire [72:0] between_9_1;
wire [72:0] between_10_1;
wire [72:0] between_11_1;
wire [72:0] between_12_1;
wire [72:0] between_13_1;
wire [72:0] between_14_1;
wire [72:0] between_15_1;
wire [72:0] between_0_2;
wire [72:0] between_1_2;
wire [72:0] between_2_2;
wire [72:0] between_3_2;
wire [72:0] between_4_2;
wire [72:0] between_5_2;
wire [72:0] between_6_2;
wire [72:0] between_7_2;
wire [72:0] between_8_2;
wire [72:0] between_9_2;
wire [72:0] between_10_2;
wire [72:0] between_11_2;
wire [72:0] between_12_2;
wire [72:0] between_13_2;
wire [72:0] between_14_2;
wire [72:0] between_15_2;
wire [72:0] between_0_3;
wire [72:0] between_1_3;
wire [72:0] between_2_3;
wire [72:0] between_3_3;
wire [72:0] between_4_3;
wire [72:0] between_5_3;
wire [72:0] between_6_3;
wire [72:0] between_7_3;
wire [72:0] between_8_3;
wire [72:0] between_9_3;
wire [72:0] between_10_3;
wire [72:0] between_11_3;
wire [72:0] between_12_3;
wire [72:0] between_13_3;
wire [72:0] between_14_3;
wire [72:0] between_15_3;
reg [72:0] between_0_0_reg = 0;
reg [72:0] between_1_0_reg = 0;
reg [72:0] between_2_0_reg = 0;
reg [72:0] between_3_0_reg = 0;
reg [72:0] between_4_0_reg = 0;
reg [72:0] between_5_0_reg = 0;
reg [72:0] between_6_0_reg = 0;
reg [72:0] between_7_0_reg = 0;
reg [72:0] between_8_0_reg = 0;
reg [72:0] between_9_0_reg = 0;
reg [72:0] between_10_0_reg = 0;
reg [72:0] between_11_0_reg = 0;
reg [72:0] between_12_0_reg = 0;
reg [72:0] between_13_0_reg = 0;
reg [72:0] between_14_0_reg = 0;
reg [72:0] between_15_0_reg = 0;
reg [72:0] between_0_1_reg = 0;
reg [72:0] between_1_1_reg = 0;
reg [72:0] between_2_1_reg = 0;
reg [72:0] between_3_1_reg = 0;
reg [72:0] between_4_1_reg = 0;
reg [72:0] between_5_1_reg = 0;
reg [72:0] between_6_1_reg = 0;
reg [72:0] between_7_1_reg = 0;
reg [72:0] between_8_1_reg = 0;
reg [72:0] between_9_1_reg = 0;
reg [72:0] between_10_1_reg = 0;
reg [72:0] between_11_1_reg = 0;
reg [72:0] between_12_1_reg = 0;
reg [72:0] between_13_1_reg = 0;
reg [72:0] between_14_1_reg = 0;
reg [72:0] between_15_1_reg = 0;
reg [72:0] between_0_2_reg = 0;
reg [72:0] between_1_2_reg = 0;
reg [72:0] between_2_2_reg = 0;
reg [72:0] between_3_2_reg = 0;
reg [72:0] between_4_2_reg = 0;
reg [72:0] between_5_2_reg = 0;
reg [72:0] between_6_2_reg = 0;
reg [72:0] between_7_2_reg = 0;
reg [72:0] between_8_2_reg = 0;
reg [72:0] between_9_2_reg = 0;
reg [72:0] between_10_2_reg = 0;
reg [72:0] between_11_2_reg = 0;
reg [72:0] between_12_2_reg = 0;
reg [72:0] between_13_2_reg = 0;
reg [72:0] between_14_2_reg = 0;
reg [72:0] between_15_2_reg = 0;
reg [72:0] between_0_3_reg = 0;
reg [72:0] between_1_3_reg = 0;
reg [72:0] between_2_3_reg = 0;
reg [72:0] between_3_3_reg = 0;
reg [72:0] between_4_3_reg = 0;
reg [72:0] between_5_3_reg = 0;
reg [72:0] between_6_3_reg = 0;
reg [72:0] between_7_3_reg = 0;
reg [72:0] between_8_3_reg = 0;
reg [72:0] between_9_3_reg = 0;
reg [72:0] between_10_3_reg = 0;
reg [72:0] between_11_3_reg = 0;
reg [72:0] between_12_3_reg = 0;
reg [72:0] between_13_3_reg = 0;
reg [72:0] between_14_3_reg = 0;
reg [72:0] between_15_3_reg = 0;
/*verilator lint_off WIDTH*/
/*verilator tracing_off*/
TNT_BIN_HC0_JaSJ17_68_16_0 TNT_BIN_HC0_JaSJ17_68_16_0_instance (.in0(internal_in0), .in1(internal_in1), .in2(internal_in2), .in3(internal_in3), .in4(internal_in4), .in5(internal_in5), .in6(internal_in6), .in7(internal_in7), .in8(internal_in8), .in9(internal_in9), .in10(internal_in10), .in11(internal_in11), .in12(internal_in12), .in13(internal_in13), .in14(internal_in14), .in15(internal_in15), .out0(between_0_0), .out1(between_1_0), .out2(between_2_0), .out3(between_3_0), .out4(between_4_0), .out5(between_5_0), .out6(between_6_0), .out7(between_7_0), .out8(between_8_0), .out9(between_9_0), .out10(between_10_0), .out11(between_11_0), .out12(between_12_0), .out13(between_13_0), .out14(between_14_0), .out15(between_15_0));
TNT_BIN_HC0_JaSJ17_68_16_1 TNT_BIN_HC0_JaSJ17_68_16_1_instance (.in0(between_0_0_reg), .in1(between_1_0_reg), .in2(between_2_0_reg), .in3(between_3_0_reg), .in4(between_4_0_reg), .in5(between_5_0_reg), .in6(between_6_0_reg), .in7(between_7_0_reg), .in8(between_8_0_reg), .in9(between_9_0_reg), .in10(between_10_0_reg), .in11(between_11_0_reg), .in12(between_12_0_reg), .in13(between_13_0_reg), .in14(between_14_0_reg), .in15(between_15_0_reg), .out0(between_0_1), .out1(between_1_1), .out2(between_2_1), .out3(between_3_1), .out4(between_4_1), .out5(between_5_1), .out6(between_6_1), .out7(between_7_1), .out8(between_8_1), .out9(between_9_1), .out10(between_10_1), .out11(between_11_1), .out12(between_12_1), .out13(between_13_1), .out14(between_14_1), .out15(between_15_1));
TNT_BIN_HC0_JaSJ17_68_16_2 TNT_BIN_HC0_JaSJ17_68_16_2_instance (.in0(between_0_1_reg), .in1(between_1_1_reg), .in2(between_2_1_reg), .in3(between_3_1_reg), .in4(between_4_1_reg), .in5(between_5_1_reg), .in6(between_6_1_reg), .in7(between_7_1_reg), .in8(between_8_1_reg), .in9(between_9_1_reg), .in10(between_10_1_reg), .in11(between_11_1_reg), .in12(between_12_1_reg), .in13(between_13_1_reg), .in14(between_14_1_reg), .in15(between_15_1_reg), .out0(between_0_2), .out1(between_1_2), .out2(between_2_2), .out3(between_3_2), .out4(between_4_2), .out5(between_5_2), .out6(between_6_2), .out7(between_7_2), .out8(between_8_2), .out9(between_9_2), .out10(between_10_2), .out11(between_11_2), .out12(between_12_2), .out13(between_13_2), .out14(between_14_2), .out15(between_15_2));
TNT_BIN_HC0_JaSJ17_68_16_3 TNT_BIN_HC0_JaSJ17_68_16_3_instance (.in0(between_0_2_reg), .in1(between_1_2_reg), .in2(between_2_2_reg), .in3(between_3_2_reg), .in4(between_4_2_reg), .in5(between_5_2_reg), .in6(between_6_2_reg), .in7(between_7_2_reg), .in8(between_8_2_reg), .in9(between_9_2_reg), .in10(between_10_2_reg), .in11(between_11_2_reg), .in12(between_12_2_reg), .in13(between_13_2_reg), .in14(between_14_2_reg), .in15(between_15_2_reg), .out0(between_0_3), .out1(between_1_3), .out2(between_2_3), .out3(between_3_3), .out4(between_4_3), .out5(between_5_3), .out6(between_6_3), .out7(between_7_3), .out8(between_8_3), .out9(between_9_3), .out10(between_10_3), .out11(between_11_3), .out12(between_12_3), .out13(between_13_3), .out14(between_14_3), .out15(between_15_3));
TNT_BIN_HC0_JaSJ17_68_16_4 TNT_BIN_HC0_JaSJ17_68_16_4_instance (.in0(between_0_3_reg), .in1(between_1_3_reg), .in2(between_2_3_reg), .in3(between_3_3_reg), .in4(between_4_3_reg), .in5(between_5_3_reg), .in6(between_6_3_reg), .in7(between_7_3_reg), .in8(between_8_3_reg), .in9(between_9_3_reg), .in10(between_10_3_reg), .in11(between_11_3_reg), .in12(between_12_3_reg), .in13(between_13_3_reg), .in14(between_14_3_reg), .in15(between_15_3_reg), .out0(internal_out0), .out1(internal_out1), .out2(internal_out2), .out3(internal_out3), .out4(internal_out4), .out5(internal_out5), .out6(internal_out6), .out7(internal_out7), .out8(internal_out8), .out9(internal_out9), .out10(internal_out10), .out11(internal_out11), .out12(internal_out12), .out13(internal_out13), .out14(internal_out14), .out15(internal_out15));
/*verilator tracing_on*/
/*verilator lint_on WIDTH*/
assign out0.from = internal_out0[67:64];
assign out0.to = 0;
assign out0.data = internal_out0[63:0];
assign out0.valid = internal_out0[68];
assign out1.from = internal_out1[67:64];
assign out1.to = 1;
assign out1.data = internal_out1[63:0];
assign out1.valid = internal_out1[68];
assign out2.from = internal_out2[67:64];
assign out2.to = 2;
assign out2.data = internal_out2[63:0];
assign out2.valid = internal_out2[68];
assign out3.from = internal_out3[67:64];
assign out3.to = 3;
assign out3.data = internal_out3[63:0];
assign out3.valid = internal_out3[68];
assign out4.from = internal_out4[67:64];
assign out4.to = 4;
assign out4.data = internal_out4[63:0];
assign out4.valid = internal_out4[68];
assign out5.from = internal_out5[67:64];
assign out5.to = 5;
assign out5.data = internal_out5[63:0];
assign out5.valid = internal_out5[68];
assign out6.from = internal_out6[67:64];
assign out6.to = 6;
assign out6.data = internal_out6[63:0];
assign out6.valid = internal_out6[68];
assign out7.from = internal_out7[67:64];
assign out7.to = 7;
assign out7.data = internal_out7[63:0];
assign out7.valid = internal_out7[68];
assign out8.from = internal_out8[67:64];
assign out8.to = 8;
assign out8.data = internal_out8[63:0];
assign out8.valid = internal_out8[68];
assign out9.from = internal_out9[67:64];
assign out9.to = 9;
assign out9.data = internal_out9[63:0];
assign out9.valid = internal_out9[68];
assign out10.from = internal_out10[67:64];
assign out10.to = 10;
assign out10.data = internal_out10[63:0];
assign out10.valid = internal_out10[68];
assign out11.from = internal_out11[67:64];
assign out11.to = 11;
assign out11.data = internal_out11[63:0];
assign out11.valid = internal_out11[68];
assign out12.from = internal_out12[67:64];
assign out12.to = 12;
assign out12.data = internal_out12[63:0];
assign out12.valid = internal_out12[68];
assign out13.from = internal_out13[67:64];
assign out13.to = 13;
assign out13.data = internal_out13[63:0];
assign out13.valid = internal_out13[68];
assign out14.from = internal_out14[67:64];
assign out14.to = 14;
assign out14.data = internal_out14[63:0];
assign out14.valid = internal_out14[68];
assign out15.from = internal_out15[67:64];
assign out15.to = 15;
assign out15.data = internal_out15[63:0];
assign out15.valid = internal_out15[68];
assign internal_in0[67:64] = in0.from;
assign internal_in0[72:69] = in0.to;
assign internal_in0[63:0] = in0.data;
assign internal_in0[68] = in0.valid;
assign internal_in1[67:64] = in1.from;
assign internal_in1[72:69] = in1.to;
assign internal_in1[63:0] = in1.data;
assign internal_in1[68] = in1.valid;
assign internal_in2[67:64] = in2.from;
assign internal_in2[72:69] = in2.to;
assign internal_in2[63:0] = in2.data;
assign internal_in2[68] = in2.valid;
assign internal_in3[67:64] = in3.from;
assign internal_in3[72:69] = in3.to;
assign internal_in3[63:0] = in3.data;
assign internal_in3[68] = in3.valid;
assign internal_in4[67:64] = in4.from;
assign internal_in4[72:69] = in4.to;
assign internal_in4[63:0] = in4.data;
assign internal_in4[68] = in4.valid;
assign internal_in5[67:64] = in5.from;
assign internal_in5[72:69] = in5.to;
assign internal_in5[63:0] = in5.data;
assign internal_in5[68] = in5.valid;
assign internal_in6[67:64] = in6.from;
assign internal_in6[72:69] = in6.to;
assign internal_in6[63:0] = in6.data;
assign internal_in6[68] = in6.valid;
assign internal_in7[67:64] = in7.from;
assign internal_in7[72:69] = in7.to;
assign internal_in7[63:0] = in7.data;
assign internal_in7[68] = in7.valid;
assign internal_in8[67:64] = in8.from;
assign internal_in8[72:69] = in8.to;
assign internal_in8[63:0] = in8.data;
assign internal_in8[68] = in8.valid;
assign internal_in9[67:64] = in9.from;
assign internal_in9[72:69] = in9.to;
assign internal_in9[63:0] = in9.data;
assign internal_in9[68] = in9.valid;
assign internal_in10[67:64] = in10.from;
assign internal_in10[72:69] = in10.to;
assign internal_in10[63:0] = in10.data;
assign internal_in10[68] = in10.valid;
assign internal_in11[67:64] = in11.from;
assign internal_in11[72:69] = in11.to;
assign internal_in11[63:0] = in11.data;
assign internal_in11[68] = in11.valid;
assign internal_in12[67:64] = in12.from;
assign internal_in12[72:69] = in12.to;
assign internal_in12[63:0] = in12.data;
assign internal_in12[68] = in12.valid;
assign internal_in13[67:64] = in13.from;
assign internal_in13[72:69] = in13.to;
assign internal_in13[63:0] = in13.data;
assign internal_in13[68] = in13.valid;
assign internal_in14[67:64] = in14.from;
assign internal_in14[72:69] = in14.to;
assign internal_in14[63:0] = in14.data;
assign internal_in14[68] = in14.valid;
assign internal_in15[67:64] = in15.from;
assign internal_in15[72:69] = in15.to;
assign internal_in15[63:0] = in15.data;
assign internal_in15[68] = in15.valid;
always @ (posedge clock) begin
  between_0_0_reg <= between_0_0;
  between_1_0_reg <= between_1_0;
  between_2_0_reg <= between_2_0;
  between_3_0_reg <= between_3_0;
  between_4_0_reg <= between_4_0;
  between_5_0_reg <= between_5_0;
  between_6_0_reg <= between_6_0;
  between_7_0_reg <= between_7_0;
  between_8_0_reg <= between_8_0;
  between_9_0_reg <= between_9_0;
  between_10_0_reg <= between_10_0;
  between_11_0_reg <= between_11_0;
  between_12_0_reg <= between_12_0;
  between_13_0_reg <= between_13_0;
  between_14_0_reg <= between_14_0;
  between_15_0_reg <= between_15_0;
  between_0_1_reg <= between_0_1;
  between_1_1_reg <= between_1_1;
  between_2_1_reg <= between_2_1;
  between_3_1_reg <= between_3_1;
  between_4_1_reg <= between_4_1;
  between_5_1_reg <= between_5_1;
  between_6_1_reg <= between_6_1;
  between_7_1_reg <= between_7_1;
  between_8_1_reg <= between_8_1;
  between_9_1_reg <= between_9_1;
  between_10_1_reg <= between_10_1;
  between_11_1_reg <= between_11_1;
  between_12_1_reg <= between_12_1;
  between_13_1_reg <= between_13_1;
  between_14_1_reg <= between_14_1;
  between_15_1_reg <= between_15_1;
  between_0_2_reg <= between_0_2;
  between_1_2_reg <= between_1_2;
  between_2_2_reg <= between_2_2;
  between_3_2_reg <= between_3_2;
  between_4_2_reg <= between_4_2;
  between_5_2_reg <= between_5_2;
  between_6_2_reg <= between_6_2;
  between_7_2_reg <= between_7_2;
  between_8_2_reg <= between_8_2;
  between_9_2_reg <= between_9_2;
  between_10_2_reg <= between_10_2;
  between_11_2_reg <= between_11_2;
  between_12_2_reg <= between_12_2;
  between_13_2_reg <= between_13_2;
  between_14_2_reg <= between_14_2;
  between_15_2_reg <= between_15_2;
  between_0_3_reg <= between_0_3;
  between_1_3_reg <= between_1_3;
  between_2_3_reg <= between_2_3;
  between_3_3_reg <= between_3_3;
  between_4_3_reg <= between_4_3;
  between_5_3_reg <= between_5_3;
  between_6_3_reg <= between_6_3;
  between_7_3_reg <= between_7_3;
  between_8_3_reg <= between_8_3;
  between_9_3_reg <= between_9_3;
  between_10_3_reg <= between_10_3;
  between_11_3_reg <= between_11_3;
  between_12_3_reg <= between_12_3;
  between_13_3_reg <= between_13_3;
  between_14_3_reg <= between_14_3;
  between_15_3_reg <= between_15_3;
end
`ifdef FORMAL
unique_destination: assume property ((!(in0.valid && in1.valid) || (in0.to != in1.to)) && (!(in0.valid && in2.valid) || (in0.to != in2.to)) && (!(in0.valid && in3.valid) || (in0.to != in3.to)) && (!(in0.valid && in4.valid) || (in0.to != in4.to)) && (!(in0.valid && in5.valid) || (in0.to != in5.to)) && (!(in0.valid && in6.valid) || (in0.to != in6.to)) && (!(in0.valid && in7.valid) || (in0.to != in7.to)) && (!(in0.valid && in8.valid) || (in0.to != in8.to)) && (!(in0.valid && in9.valid) || (in0.to != in9.to)) && (!(in0.valid && in10.valid) || (in0.to != in10.to)) && (!(in0.valid && in11.valid) || (in0.to != in11.to)) && (!(in0.valid && in12.valid) || (in0.to != in12.to)) && (!(in0.valid && in13.valid) || (in0.to != in13.to)) && (!(in0.valid && in14.valid) || (in0.to != in14.to)) && (!(in0.valid && in15.valid) || (in0.to != in15.to)) && (!(in1.valid && in0.valid) || (in1.to != in0.to)) && (!(in1.valid && in2.valid) || (in1.to != in2.to)) && (!(in1.valid && in3.valid) || (in1.to != in3.to)) && (!(in1.valid && in4.valid) || (in1.to != in4.to)) && (!(in1.valid && in5.valid) || (in1.to != in5.to)) && (!(in1.valid && in6.valid) || (in1.to != in6.to)) && (!(in1.valid && in7.valid) || (in1.to != in7.to)) && (!(in1.valid && in8.valid) || (in1.to != in8.to)) && (!(in1.valid && in9.valid) || (in1.to != in9.to)) && (!(in1.valid && in10.valid) || (in1.to != in10.to)) && (!(in1.valid && in11.valid) || (in1.to != in11.to)) && (!(in1.valid && in12.valid) || (in1.to != in12.to)) && (!(in1.valid && in13.valid) || (in1.to != in13.to)) && (!(in1.valid && in14.valid) || (in1.to != in14.to)) && (!(in1.valid && in15.valid) || (in1.to != in15.to)) && (!(in2.valid && in0.valid) || (in2.to != in0.to)) && (!(in2.valid && in1.valid) || (in2.to != in1.to)) && (!(in2.valid && in3.valid) || (in2.to != in3.to)) && (!(in2.valid && in4.valid) || (in2.to != in4.to)) && (!(in2.valid && in5.valid) || (in2.to != in5.to)) && (!(in2.valid && in6.valid) || (in2.to != in6.to)) && (!(in2.valid && in7.valid) || (in2.to != in7.to)) && (!(in2.valid && in8.valid) || (in2.to != in8.to)) && (!(in2.valid && in9.valid) || (in2.to != in9.to)) && (!(in2.valid && in10.valid) || (in2.to != in10.to)) && (!(in2.valid && in11.valid) || (in2.to != in11.to)) && (!(in2.valid && in12.valid) || (in2.to != in12.to)) && (!(in2.valid && in13.valid) || (in2.to != in13.to)) && (!(in2.valid && in14.valid) || (in2.to != in14.to)) && (!(in2.valid && in15.valid) || (in2.to != in15.to)) && (!(in3.valid && in0.valid) || (in3.to != in0.to)) && (!(in3.valid && in1.valid) || (in3.to != in1.to)) && (!(in3.valid && in2.valid) || (in3.to != in2.to)) && (!(in3.valid && in4.valid) || (in3.to != in4.to)) && (!(in3.valid && in5.valid) || (in3.to != in5.to)) && (!(in3.valid && in6.valid) || (in3.to != in6.to)) && (!(in3.valid && in7.valid) || (in3.to != in7.to)) && (!(in3.valid && in8.valid) || (in3.to != in8.to)) && (!(in3.valid && in9.valid) || (in3.to != in9.to)) && (!(in3.valid && in10.valid) || (in3.to != in10.to)) && (!(in3.valid && in11.valid) || (in3.to != in11.to)) && (!(in3.valid && in12.valid) || (in3.to != in12.to)) && (!(in3.valid && in13.valid) || (in3.to != in13.to)) && (!(in3.valid && in14.valid) || (in3.to != in14.to)) && (!(in3.valid && in15.valid) || (in3.to != in15.to)) && (!(in4.valid && in0.valid) || (in4.to != in0.to)) && (!(in4.valid && in1.valid) || (in4.to != in1.to)) && (!(in4.valid && in2.valid) || (in4.to != in2.to)) && (!(in4.valid && in3.valid) || (in4.to != in3.to)) && (!(in4.valid && in5.valid) || (in4.to != in5.to)) && (!(in4.valid && in6.valid) || (in4.to != in6.to)) && (!(in4.valid && in7.valid) || (in4.to != in7.to)) && (!(in4.valid && in8.valid) || (in4.to != in8.to)) && (!(in4.valid && in9.valid) || (in4.to != in9.to)) && (!(in4.valid && in10.valid) || (in4.to != in10.to)) && (!(in4.valid && in11.valid) || (in4.to != in11.to)) && (!(in4.valid && in12.valid) || (in4.to != in12.to)) && (!(in4.valid && in13.valid) || (in4.to != in13.to)) && (!(in4.valid && in14.valid) || (in4.to != in14.to)) && (!(in4.valid && in15.valid) || (in4.to != in15.to)) && (!(in5.valid && in0.valid) || (in5.to != in0.to)) && (!(in5.valid && in1.valid) || (in5.to != in1.to)) && (!(in5.valid && in2.valid) || (in5.to != in2.to)) && (!(in5.valid && in3.valid) || (in5.to != in3.to)) && (!(in5.valid && in4.valid) || (in5.to != in4.to)) && (!(in5.valid && in6.valid) || (in5.to != in6.to)) && (!(in5.valid && in7.valid) || (in5.to != in7.to)) && (!(in5.valid && in8.valid) || (in5.to != in8.to)) && (!(in5.valid && in9.valid) || (in5.to != in9.to)) && (!(in5.valid && in10.valid) || (in5.to != in10.to)) && (!(in5.valid && in11.valid) || (in5.to != in11.to)) && (!(in5.valid && in12.valid) || (in5.to != in12.to)) && (!(in5.valid && in13.valid) || (in5.to != in13.to)) && (!(in5.valid && in14.valid) || (in5.to != in14.to)) && (!(in5.valid && in15.valid) || (in5.to != in15.to)) && (!(in6.valid && in0.valid) || (in6.to != in0.to)) && (!(in6.valid && in1.valid) || (in6.to != in1.to)) && (!(in6.valid && in2.valid) || (in6.to != in2.to)) && (!(in6.valid && in3.valid) || (in6.to != in3.to)) && (!(in6.valid && in4.valid) || (in6.to != in4.to)) && (!(in6.valid && in5.valid) || (in6.to != in5.to)) && (!(in6.valid && in7.valid) || (in6.to != in7.to)) && (!(in6.valid && in8.valid) || (in6.to != in8.to)) && (!(in6.valid && in9.valid) || (in6.to != in9.to)) && (!(in6.valid && in10.valid) || (in6.to != in10.to)) && (!(in6.valid && in11.valid) || (in6.to != in11.to)) && (!(in6.valid && in12.valid) || (in6.to != in12.to)) && (!(in6.valid && in13.valid) || (in6.to != in13.to)) && (!(in6.valid && in14.valid) || (in6.to != in14.to)) && (!(in6.valid && in15.valid) || (in6.to != in15.to)) && (!(in7.valid && in0.valid) || (in7.to != in0.to)) && (!(in7.valid && in1.valid) || (in7.to != in1.to)) && (!(in7.valid && in2.valid) || (in7.to != in2.to)) && (!(in7.valid && in3.valid) || (in7.to != in3.to)) && (!(in7.valid && in4.valid) || (in7.to != in4.to)) && (!(in7.valid && in5.valid) || (in7.to != in5.to)) && (!(in7.valid && in6.valid) || (in7.to != in6.to)) && (!(in7.valid && in8.valid) || (in7.to != in8.to)) && (!(in7.valid && in9.valid) || (in7.to != in9.to)) && (!(in7.valid && in10.valid) || (in7.to != in10.to)) && (!(in7.valid && in11.valid) || (in7.to != in11.to)) && (!(in7.valid && in12.valid) || (in7.to != in12.to)) && (!(in7.valid && in13.valid) || (in7.to != in13.to)) && (!(in7.valid && in14.valid) || (in7.to != in14.to)) && (!(in7.valid && in15.valid) || (in7.to != in15.to)) && (!(in8.valid && in0.valid) || (in8.to != in0.to)) && (!(in8.valid && in1.valid) || (in8.to != in1.to)) && (!(in8.valid && in2.valid) || (in8.to != in2.to)) && (!(in8.valid && in3.valid) || (in8.to != in3.to)) && (!(in8.valid && in4.valid) || (in8.to != in4.to)) && (!(in8.valid && in5.valid) || (in8.to != in5.to)) && (!(in8.valid && in6.valid) || (in8.to != in6.to)) && (!(in8.valid && in7.valid) || (in8.to != in7.to))
        && (!(in8.valid && in9.valid) || (in8.to != in9.to)) && (!(in8.valid && in10.valid) || (in8.to != in10.to)) && (!(in8.valid && in11.valid) || (in8.to != in11.to)) && (!(in8.valid && in12.valid) || (in8.to != in12.to)) && (!(in8.valid && in13.valid) || (in8.to != in13.to)) && (!(in8.valid && in14.valid) || (in8.to != in14.to)) && (!(in8.valid && in15.valid) || (in8.to != in15.to)) && (!(in9.valid && in0.valid) || (in9.to != in0.to)) && (!(in9.valid && in1.valid) || (in9.to != in1.to)) && (!(in9.valid && in2.valid) || (in9.to != in2.to)) && (!(in9.valid && in3.valid) || (in9.to != in3.to)) && (!(in9.valid && in4.valid) || (in9.to != in4.to)) && (!(in9.valid && in5.valid) || (in9.to != in5.to)) && (!(in9.valid && in6.valid) || (in9.to != in6.to)) && (!(in9.valid && in7.valid) || (in9.to != in7.to)) && (!(in9.valid && in8.valid) || (in9.to != in8.to)) && (!(in9.valid && in10.valid) || (in9.to != in10.to)) && (!(in9.valid && in11.valid) || (in9.to != in11.to)) && (!(in9.valid && in12.valid) || (in9.to != in12.to)) && (!(in9.valid && in13.valid) || (in9.to != in13.to)) && (!(in9.valid && in14.valid) || (in9.to != in14.to)) && (!(in9.valid && in15.valid) || (in9.to != in15.to)) && (!(in10.valid && in0.valid) || (in10.to != in0.to)) && (!(in10.valid && in1.valid) || (in10.to != in1.to)) && (!(in10.valid && in2.valid) || (in10.to != in2.to)) && (!(in10.valid && in3.valid) || (in10.to != in3.to)) && (!(in10.valid && in4.valid) || (in10.to != in4.to)) && (!(in10.valid && in5.valid) || (in10.to != in5.to)) && (!(in10.valid && in6.valid) || (in10.to != in6.to)) && (!(in10.valid && in7.valid) || (in10.to != in7.to)) && (!(in10.valid && in8.valid) || (in10.to != in8.to)) && (!(in10.valid && in9.valid) || (in10.to != in9.to)) && (!(in10.valid && in11.valid) || (in10.to != in11.to)) && (!(in10.valid && in12.valid) || (in10.to != in12.to)) && (!(in10.valid && in13.valid) || (in10.to != in13.to)) && (!(in10.valid && in14.valid) || (in10.to != in14.to)) && (!(in10.valid && in15.valid) || (in10.to != in15.to)) && (!(in11.valid && in0.valid) || (in11.to != in0.to)) && (!(in11.valid && in1.valid) || (in11.to != in1.to)) && (!(in11.valid && in2.valid) || (in11.to != in2.to)) && (!(in11.valid && in3.valid) || (in11.to != in3.to)) && (!(in11.valid && in4.valid) || (in11.to != in4.to)) && (!(in11.valid && in5.valid) || (in11.to != in5.to)) && (!(in11.valid && in6.valid) || (in11.to != in6.to)) && (!(in11.valid && in7.valid) || (in11.to != in7.to)) && (!(in11.valid && in8.valid) || (in11.to != in8.to)) && (!(in11.valid && in9.valid) || (in11.to != in9.to)) && (!(in11.valid && in10.valid) || (in11.to != in10.to)) && (!(in11.valid && in12.valid) || (in11.to != in12.to)) && (!(in11.valid && in13.valid) || (in11.to != in13.to)) && (!(in11.valid && in14.valid) || (in11.to != in14.to)) && (!(in11.valid && in15.valid) || (in11.to != in15.to)) && (!(in12.valid && in0.valid) || (in12.to != in0.to)) && (!(in12.valid && in1.valid) || (in12.to != in1.to)) && (!(in12.valid && in2.valid) || (in12.to != in2.to)) && (!(in12.valid && in3.valid) || (in12.to != in3.to)) && (!(in12.valid && in4.valid) || (in12.to != in4.to)) && (!(in12.valid && in5.valid) || (in12.to != in5.to)) && (!(in12.valid && in6.valid) || (in12.to != in6.to)) && (!(in12.valid && in7.valid) || (in12.to != in7.to)) && (!(in12.valid && in8.valid) || (in12.to != in8.to)) && (!(in12.valid && in9.valid) || (in12.to != in9.to)) && (!(in12.valid && in10.valid) || (in12.to != in10.to)) && (!(in12.valid && in11.valid) || (in12.to != in11.to)) && (!(in12.valid && in13.valid) || (in12.to != in13.to)) && (!(in12.valid && in14.valid) || (in12.to != in14.to)) && (!(in12.valid && in15.valid) || (in12.to != in15.to)) && (!(in13.valid && in0.valid) || (in13.to != in0.to)) && (!(in13.valid && in1.valid) || (in13.to != in1.to)) && (!(in13.valid && in2.valid) || (in13.to != in2.to)) && (!(in13.valid && in3.valid) || (in13.to != in3.to)) && (!(in13.valid && in4.valid) || (in13.to != in4.to)) && (!(in13.valid && in5.valid) || (in13.to != in5.to)) && (!(in13.valid && in6.valid) || (in13.to != in6.to)) && (!(in13.valid && in7.valid) || (in13.to != in7.to)) && (!(in13.valid && in8.valid) || (in13.to != in8.to)) && (!(in13.valid && in9.valid) || (in13.to != in9.to)) && (!(in13.valid && in10.valid) || (in13.to != in10.to)) && (!(in13.valid && in11.valid) || (in13.to != in11.to)) && (!(in13.valid && in12.valid) || (in13.to != in12.to)) && (!(in13.valid && in14.valid) || (in13.to != in14.to)) && (!(in13.valid && in15.valid) || (in13.to != in15.to)) && (!(in14.valid && in0.valid) || (in14.to != in0.to)) && (!(in14.valid && in1.valid) || (in14.to != in1.to)) && (!(in14.valid && in2.valid) || (in14.to != in2.to)) && (!(in14.valid && in3.valid) || (in14.to != in3.to)) && (!(in14.valid && in4.valid) || (in14.to != in4.to)) && (!(in14.valid && in5.valid) || (in14.to != in5.to)) && (!(in14.valid && in6.valid) || (in14.to != in6.to)) && (!(in14.valid && in7.valid) || (in14.to != in7.to)) && (!(in14.valid && in8.valid) || (in14.to != in8.to)) && (!(in14.valid && in9.valid) || (in14.to != in9.to)) && (!(in14.valid && in10.valid) || (in14.to != in10.to)) && (!(in14.valid && in11.valid) || (in14.to != in11.to)) && (!(in14.valid && in12.valid) || (in14.to != in12.to)) && (!(in14.valid && in13.valid) || (in14.to != in13.to)) && (!(in14.valid && in15.valid) || (in14.to != in15.to)) && (!(in15.valid && in0.valid) || (in15.to != in0.to)) && (!(in15.valid && in1.valid) || (in15.to != in1.to)) && (!(in15.valid && in2.valid) || (in15.to != in2.to)) && (!(in15.valid && in3.valid) || (in15.to != in3.to)) && (!(in15.valid && in4.valid) || (in15.to != in4.to)) && (!(in15.valid && in5.valid) || (in15.to != in5.to)) && (!(in15.valid && in6.valid) || (in15.to != in6.to)) && (!(in15.valid && in7.valid) || (in15.to != in7.to)) && (!(in15.valid && in8.valid) || (in15.to != in8.to)) && (!(in15.valid && in9.valid) || (in15.to != in9.to)) && (!(in15.valid && in10.valid) || (in15.to != in10.to)) && (!(in15.valid && in11.valid) || (in15.to != in11.to)) && (!(in15.valid && in12.valid) || (in15.to != in12.to)) && (!(in15.valid && in13.valid) || (in15.to != in13.to)) && (!(in15.valid && in14.valid) || (in15.to != in14.to)));
correct_from: assume property ((!in0.valid || (in0.from == 0)) && (!in1.valid || (in1.from == 1)) && (!in2.valid || (in2.from == 2)) && (!in3.valid || (in3.from == 3)) && (!in4.valid || (in4.from == 4)) && (!in5.valid || (in5.from == 5)) && (!in6.valid || (in6.from == 6)) && (!in7.valid || (in7.from == 7)) && (!in8.valid || (in8.from == 8)) && (!in9.valid || (in9.from == 9)) && (!in10.valid || (in10.from == 10)) && (!in11.valid || (in11.from == 11)) && (!in12.valid || (in12.from == 12)) && (!in13.valid || (in13.from == 13)) && (!in14.valid || (in14.from == 14)) && (!in15.valid || (in15.from == 15)));
correct_dest: assume property ((!in0.valid || (in0.to < 16)) && (!in1.valid || (in1.to < 16)) && (!in2.valid || (in2.to < 16)) && (!in3.valid || (in3.to < 16)) && (!in4.valid || (in4.to < 16)) && (!in5.valid || (in5.to < 16)) && (!in6.valid || (in6.to < 16)) && (!in7.valid || (in7.to < 16)) && (!in8.valid || (in8.to < 16)) && (!in9.valid || (in9.to < 16)) && (!in10.valid || (in10.to < 16)) && (!in11.valid || (in11.to < 16)) && (!in12.valid || (in12.to < 16)) && (!in13.valid || (in13.to < 16)) && (!in14.valid || (in14.to < 16)) && (!in15.valid || (in15.to < 16)));
reg [$clog2(5)-1:0] proof_cycles = 0;
always @ (posedge clock) begin
  if (proof_cycles < 4) begin
    proof_cycles <= proof_cycles + 1;
    all_ports_starting_invalid: assert (!out0.valid && !out1.valid && !out2.valid && !out3.valid && !out4.valid && !out5.valid && !out6.valid && !out7.valid && !out8.valid && !out9.valid && !out10.valid && !out11.valid && !out12.valid && !out13.valid && !out14.valid && !out15.valid);
  end else begin
    // Sanity checks.
    all_outputs_valid: cover (out0.valid && out1.valid && out2.valid && out3.valid && out4.valid && out5.valid && out6.valid && out7.valid && out8.valid && out9.valid && out10.valid && out11.valid && out12.valid && out13.valid && out14.valid && out15.valid);
    // Goals of implementation.
    correct_source_exists: assert ((!out0.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 0) && ($past(in0.data, 4) == out0.data) && (out0.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 0) && ($past(in1.data, 4) == out0.data) && (out0.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 0) && ($past(in2.data, 4) == out0.data) && (out0.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 0) && ($past(in3.data, 4) == out0.data) && (out0.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 0) && ($past(in4.data, 4) == out0.data) && (out0.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 0) && ($past(in5.data, 4) == out0.data) && (out0.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 0) && ($past(in6.data, 4) == out0.data) && (out0.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 0) && ($past(in7.data, 4) == out0.data) && (out0.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 0) && ($past(in8.data, 4) == out0.data) && (out0.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 0) && ($past(in9.data, 4) == out0.data) && (out0.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 0) && ($past(in10.data, 4) == out0.data) && (out0.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 0) && ($past(in11.data, 4) == out0.data) && (out0.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 0) && ($past(in12.data, 4) == out0.data) && (out0.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 0) && ($past(in13.data, 4) == out0.data) && (out0.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 0) && ($past(in14.data, 4) == out0.data) && (out0.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 0) && ($past(in15.data, 4) == out0.data) && (out0.from == 15))))
        && (!out1.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 1) && ($past(in0.data, 4) == out1.data) && (out1.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 1) && ($past(in1.data, 4) == out1.data) && (out1.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 1) && ($past(in2.data, 4) == out1.data) && (out1.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 1) && ($past(in3.data, 4) == out1.data) && (out1.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 1) && ($past(in4.data, 4) == out1.data) && (out1.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 1) && ($past(in5.data, 4) == out1.data) && (out1.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 1) && ($past(in6.data, 4) == out1.data) && (out1.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 1) && ($past(in7.data, 4) == out1.data) && (out1.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 1) && ($past(in8.data, 4) == out1.data) && (out1.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 1) && ($past(in9.data, 4) == out1.data) && (out1.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 1) && ($past(in10.data, 4) == out1.data) && (out1.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 1) && ($past(in11.data, 4) == out1.data) && (out1.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 1) && ($past(in12.data, 4) == out1.data) && (out1.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 1) && ($past(in13.data, 4) == out1.data) && (out1.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 1) && ($past(in14.data, 4) == out1.data) && (out1.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 1) && ($past(in15.data, 4) == out1.data) && (out1.from == 15))))
        && (!out2.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 2) && ($past(in0.data, 4) == out2.data) && (out2.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 2) && ($past(in1.data, 4) == out2.data) && (out2.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 2) && ($past(in2.data, 4) == out2.data) && (out2.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 2) && ($past(in3.data, 4) == out2.data) && (out2.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 2) && ($past(in4.data, 4) == out2.data) && (out2.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 2) && ($past(in5.data, 4) == out2.data) && (out2.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 2) && ($past(in6.data, 4) == out2.data) && (out2.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 2) && ($past(in7.data, 4) == out2.data) && (out2.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 2) && ($past(in8.data, 4) == out2.data) && (out2.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 2) && ($past(in9.data, 4) == out2.data) && (out2.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 2) && ($past(in10.data, 4) == out2.data) && (out2.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 2) && ($past(in11.data, 4) == out2.data) && (out2.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 2) && ($past(in12.data, 4) == out2.data) && (out2.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 2) && ($past(in13.data, 4) == out2.data) && (out2.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 2) && ($past(in14.data, 4) == out2.data) && (out2.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 2) && ($past(in15.data, 4) == out2.data) && (out2.from == 15))))
        && (!out3.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 3) && ($past(in0.data, 4) == out3.data) && (out3.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 3) && ($past(in1.data, 4) == out3.data) && (out3.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 3) && ($past(in2.data, 4) == out3.data) && (out3.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 3) && ($past(in3.data, 4) == out3.data) && (out3.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 3) && ($past(in4.data, 4) == out3.data) && (out3.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 3) && ($past(in5.data, 4) == out3.data) && (out3.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 3) && ($past(in6.data, 4) == out3.data) && (out3.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 3) && ($past(in7.data, 4) == out3.data) && (out3.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 3) && ($past(in8.data, 4) == out3.data) && (out3.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 3) && ($past(in9.data, 4) == out3.data) && (out3.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 3) && ($past(in10.data, 4) == out3.data) && (out3.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 3) && ($past(in11.data, 4) == out3.data) && (out3.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 3) && ($past(in12.data, 4) == out3.data) && (out3.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 3) && ($past(in13.data, 4) == out3.data) && (out3.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 3) && ($past(in14.data, 4) == out3.data) && (out3.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 3) && ($past(in15.data, 4) == out3.data) && (out3.from == 15))))
        && (!out4.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 4) && ($past(in0.data, 4) == out4.data) && (out4.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 4) && ($past(in1.data, 4) == out4.data) && (out4.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 4) && ($past(in2.data, 4) == out4.data) && (out4.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 4) && ($past(in3.data, 4) == out4.data) && (out4.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 4) && ($past(in4.data, 4) == out4.data) && (out4.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 4) && ($past(in5.data, 4) == out4.data) && (out4.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 4) && ($past(in6.data, 4) == out4.data) && (out4.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 4) && ($past(in7.data, 4) == out4.data) && (out4.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 4) && ($past(in8.data, 4) == out4.data) && (out4.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 4) && ($past(in9.data, 4) == out4.data) && (out4.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 4) && ($past(in10.data, 4) == out4.data) && (out4.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 4) && ($past(in11.data, 4) == out4.data) && (out4.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 4) && ($past(in12.data, 4) == out4.data) && (out4.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 4) && ($past(in13.data, 4) == out4.data) && (out4.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 4) && ($past(in14.data, 4) == out4.data) && (out4.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 4) && ($past(in15.data, 4) == out4.data) && (out4.from == 15))))
        && (!out5.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 5) && ($past(in0.data, 4) == out5.data) && (out5.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 5) && ($past(in1.data, 4) == out5.data) && (out5.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 5) && ($past(in2.data, 4) == out5.data) && (out5.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 5) && ($past(in3.data, 4) == out5.data) && (out5.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 5) && ($past(in4.data, 4) == out5.data) && (out5.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 5) && ($past(in5.data, 4) == out5.data) && (out5.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 5) && ($past(in6.data, 4) == out5.data) && (out5.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 5) && ($past(in7.data, 4) == out5.data) && (out5.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 5) && ($past(in8.data, 4) == out5.data) && (out5.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 5) && ($past(in9.data, 4) == out5.data) && (out5.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 5) && ($past(in10.data, 4) == out5.data) && (out5.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 5) && ($past(in11.data, 4) == out5.data) && (out5.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 5) && ($past(in12.data, 4) == out5.data) && (out5.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 5) && ($past(in13.data, 4) == out5.data) && (out5.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 5) && ($past(in14.data, 4) == out5.data) && (out5.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 5) && ($past(in15.data, 4) == out5.data) && (out5.from == 15))))
        && (!out6.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 6) && ($past(in0.data, 4) == out6.data) && (out6.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 6) && ($past(in1.data, 4) == out6.data) && (out6.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 6) && ($past(in2.data, 4) == out6.data) && (out6.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 6) && ($past(in3.data, 4) == out6.data) && (out6.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 6) && ($past(in4.data, 4) == out6.data) && (out6.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 6) && ($past(in5.data, 4) == out6.data) && (out6.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 6) && ($past(in6.data, 4) == out6.data) && (out6.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 6) && ($past(in7.data, 4) == out6.data) && (out6.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 6) && ($past(in8.data, 4) == out6.data) && (out6.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 6) && ($past(in9.data, 4) == out6.data) && (out6.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 6) && ($past(in10.data, 4) == out6.data) && (out6.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 6) && ($past(in11.data, 4) == out6.data) && (out6.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 6) && ($past(in12.data, 4) == out6.data) && (out6.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 6) && ($past(in13.data, 4) == out6.data) && (out6.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 6) && ($past(in14.data, 4) == out6.data) && (out6.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 6) && ($past(in15.data, 4) == out6.data) && (out6.from == 15))))
        && (!out7.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 7) && ($past(in0.data, 4) == out7.data) && (out7.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 7) && ($past(in1.data, 4) == out7.data) && (out7.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 7) && ($past(in2.data, 4) == out7.data) && (out7.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 7) && ($past(in3.data, 4) == out7.data) && (out7.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 7) && ($past(in4.data, 4) == out7.data) && (out7.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 7) && ($past(in5.data, 4) == out7.data) && (out7.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 7) && ($past(in6.data, 4) == out7.data) && (out7.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 7) && ($past(in7.data, 4) == out7.data) && (out7.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 7) && ($past(in8.data, 4) == out7.data) && (out7.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 7) && ($past(in9.data, 4) == out7.data) && (out7.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 7) && ($past(in10.data, 4) == out7.data) && (out7.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 7) && ($past(in11.data, 4) == out7.data) && (out7.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 7) && ($past(in12.data, 4) == out7.data) && (out7.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 7) && ($past(in13.data, 4) == out7.data) && (out7.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 7) && ($past(in14.data, 4) == out7.data) && (out7.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 7) && ($past(in15.data, 4) == out7.data) && (out7.from == 15))))
        && (!out8.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 8) && ($past(in0.data, 4) == out8.data) && (out8.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 8) && ($past(in1.data, 4) == out8.data) && (out8.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 8) && ($past(in2.data, 4) == out8.data) && (out8.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 8) && ($past(in3.data, 4) == out8.data) && (out8.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 8) && ($past(in4.data, 4) == out8.data) && (out8.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 8) && ($past(in5.data, 4) == out8.data) && (out8.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 8) && ($past(in6.data, 4) == out8.data) && (out8.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 8) && ($past(in7.data, 4) == out8.data) && (out8.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 8) && ($past(in8.data, 4) == out8.data) && (out8.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 8) && ($past(in9.data, 4) == out8.data) && (out8.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 8) && ($past(in10.data, 4) == out8.data) && (out8.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 8) && ($past(in11.data, 4) == out8.data) && (out8.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 8) && ($past(in12.data, 4) == out8.data) && (out8.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 8) && ($past(in13.data, 4) == out8.data) && (out8.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 8) && ($past(in14.data, 4) == out8.data) && (out8.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 8) && ($past(in15.data, 4) == out8.data) && (out8.from == 15))))
        && (!out9.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 9) && ($past(in0.data, 4) == out9.data) && (out9.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 9) && ($past(in1.data, 4) == out9.data) && (out9.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 9) && ($past(in2.data, 4) == out9.data) && (out9.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 9) && ($past(in3.data, 4) == out9.data) && (out9.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 9) && ($past(in4.data, 4) == out9.data) && (out9.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 9) && ($past(in5.data, 4) == out9.data) && (out9.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 9) && ($past(in6.data, 4) == out9.data) && (out9.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 9) && ($past(in7.data, 4) == out9.data) && (out9.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 9) && ($past(in8.data, 4) == out9.data) && (out9.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 9) && ($past(in9.data, 4) == out9.data) && (out9.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 9) && ($past(in10.data, 4) == out9.data) && (out9.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 9) && ($past(in11.data, 4) == out9.data) && (out9.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 9) && ($past(in12.data, 4) == out9.data) && (out9.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 9) && ($past(in13.data, 4) == out9.data) && (out9.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 9) && ($past(in14.data, 4) == out9.data) && (out9.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 9) && ($past(in15.data, 4) == out9.data) && (out9.from == 15))))
        && (!out10.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 10) && ($past(in0.data, 4) == out10.data) && (out10.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 10) && ($past(in1.data, 4) == out10.data) && (out10.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 10) && ($past(in2.data, 4) == out10.data) && (out10.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 10) && ($past(in3.data, 4) == out10.data) && (out10.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 10) && ($past(in4.data, 4) == out10.data) && (out10.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 10) && ($past(in5.data, 4) == out10.data) && (out10.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 10) && ($past(in6.data, 4) == out10.data) && (out10.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 10) && ($past(in7.data, 4) == out10.data) && (out10.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 10) && ($past(in8.data, 4) == out10.data) && (out10.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 10) && ($past(in9.data, 4) == out10.data) && (out10.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 10) && ($past(in10.data, 4) == out10.data) && (out10.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 10) && ($past(in11.data, 4) == out10.data) && (out10.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 10) && ($past(in12.data, 4) == out10.data) && (out10.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 10) && ($past(in13.data, 4) == out10.data) && (out10.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 10) && ($past(in14.data, 4) == out10.data) && (out10.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 10) && ($past(in15.data, 4) == out10.data) && (out10.from == 15))))
        && (!out11.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 11) && ($past(in0.data, 4) == out11.data) && (out11.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 11) && ($past(in1.data, 4) == out11.data) && (out11.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 11) && ($past(in2.data, 4) == out11.data) && (out11.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 11) && ($past(in3.data, 4) == out11.data) && (out11.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 11) && ($past(in4.data, 4) == out11.data) && (out11.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 11) && ($past(in5.data, 4) == out11.data) && (out11.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 11) && ($past(in6.data, 4) == out11.data) && (out11.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 11) && ($past(in7.data, 4) == out11.data) && (out11.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 11) && ($past(in8.data, 4) == out11.data) && (out11.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 11) && ($past(in9.data, 4) == out11.data) && (out11.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 11) && ($past(in10.data, 4) == out11.data) && (out11.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 11) && ($past(in11.data, 4) == out11.data) && (out11.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 11) && ($past(in12.data, 4) == out11.data) && (out11.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 11) && ($past(in13.data, 4) == out11.data) && (out11.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 11) && ($past(in14.data, 4) == out11.data) && (out11.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 11) && ($past(in15.data, 4) == out11.data) && (out11.from == 15))))
        && (!out12.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 12) && ($past(in0.data, 4) == out12.data) && (out12.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 12) && ($past(in1.data, 4) == out12.data) && (out12.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 12) && ($past(in2.data, 4) == out12.data) && (out12.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 12) && ($past(in3.data, 4) == out12.data) && (out12.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 12) && ($past(in4.data, 4) == out12.data) && (out12.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 12) && ($past(in5.data, 4) == out12.data) && (out12.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 12) && ($past(in6.data, 4) == out12.data) && (out12.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 12) && ($past(in7.data, 4) == out12.data) && (out12.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 12) && ($past(in8.data, 4) == out12.data) && (out12.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 12) && ($past(in9.data, 4) == out12.data) && (out12.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 12) && ($past(in10.data, 4) == out12.data) && (out12.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 12) && ($past(in11.data, 4) == out12.data) && (out12.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 12) && ($past(in12.data, 4) == out12.data) && (out12.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 12) && ($past(in13.data, 4) == out12.data) && (out12.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 12) && ($past(in14.data, 4) == out12.data) && (out12.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 12) && ($past(in15.data, 4) == out12.data) && (out12.from == 15))))
        && (!out13.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 13) && ($past(in0.data, 4) == out13.data) && (out13.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 13) && ($past(in1.data, 4) == out13.data) && (out13.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 13) && ($past(in2.data, 4) == out13.data) && (out13.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 13) && ($past(in3.data, 4) == out13.data) && (out13.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 13) && ($past(in4.data, 4) == out13.data) && (out13.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 13) && ($past(in5.data, 4) == out13.data) && (out13.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 13) && ($past(in6.data, 4) == out13.data) && (out13.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 13) && ($past(in7.data, 4) == out13.data) && (out13.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 13) && ($past(in8.data, 4) == out13.data) && (out13.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 13) && ($past(in9.data, 4) == out13.data) && (out13.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 13) && ($past(in10.data, 4) == out13.data) && (out13.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 13) && ($past(in11.data, 4) == out13.data) && (out13.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 13) && ($past(in12.data, 4) == out13.data) && (out13.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 13) && ($past(in13.data, 4) == out13.data) && (out13.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 13) && ($past(in14.data, 4) == out13.data) && (out13.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 13) && ($past(in15.data, 4) == out13.data) && (out13.from == 15))))
        && (!out14.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 14) && ($past(in0.data, 4) == out14.data) && (out14.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 14) && ($past(in1.data, 4) == out14.data) && (out14.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 14) && ($past(in2.data, 4) == out14.data) && (out14.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 14) && ($past(in3.data, 4) == out14.data) && (out14.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 14) && ($past(in4.data, 4) == out14.data) && (out14.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 14) && ($past(in5.data, 4) == out14.data) && (out14.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 14) && ($past(in6.data, 4) == out14.data) && (out14.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 14) && ($past(in7.data, 4) == out14.data) && (out14.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 14) && ($past(in8.data, 4) == out14.data) && (out14.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 14) && ($past(in9.data, 4) == out14.data) && (out14.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 14) && ($past(in10.data, 4) == out14.data) && (out14.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 14) && ($past(in11.data, 4) == out14.data) && (out14.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 14) && ($past(in12.data, 4) == out14.data) && (out14.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 14) && ($past(in13.data, 4) == out14.data) && (out14.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 14) && ($past(in14.data, 4) == out14.data) && (out14.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 14) && ($past(in15.data, 4) == out14.data) && (out14.from == 15))))
        && (!out15.valid || (($past(in0.valid, 4) && ($past(in0.to, 4) == 15) && ($past(in0.data, 4) == out15.data) && (out15.from == 0)) || ($past(in1.valid, 4) && ($past(in1.to, 4) == 15) && ($past(in1.data, 4) == out15.data) && (out15.from == 1)) || ($past(in2.valid, 4) && ($past(in2.to, 4) == 15) && ($past(in2.data, 4) == out15.data) && (out15.from == 2)) || ($past(in3.valid, 4) && ($past(in3.to, 4) == 15) && ($past(in3.data, 4) == out15.data) && (out15.from == 3)) || ($past(in4.valid, 4) && ($past(in4.to, 4) == 15) && ($past(in4.data, 4) == out15.data) && (out15.from == 4)) || ($past(in5.valid, 4) && ($past(in5.to, 4) == 15) && ($past(in5.data, 4) == out15.data) && (out15.from == 5)) || ($past(in6.valid, 4) && ($past(in6.to, 4) == 15) && ($past(in6.data, 4) == out15.data) && (out15.from == 6)) || ($past(in7.valid, 4) && ($past(in7.to, 4) == 15) && ($past(in7.data, 4) == out15.data) && (out15.from == 7)) || ($past(in8.valid, 4) && ($past(in8.to, 4) == 15) && ($past(in8.data, 4) == out15.data) && (out15.from == 8)) || ($past(in9.valid, 4) && ($past(in9.to, 4) == 15) && ($past(in9.data, 4) == out15.data) && (out15.from == 9)) || ($past(in10.valid, 4) && ($past(in10.to, 4) == 15) && ($past(in10.data, 4) == out15.data) && (out15.from == 10)) || ($past(in11.valid, 4) && ($past(in11.to, 4) == 15) && ($past(in11.data, 4) == out15.data) && (out15.from == 11)) || ($past(in12.valid, 4) && ($past(in12.to, 4) == 15) && ($past(in12.data, 4) == out15.data) && (out15.from == 12)) || ($past(in13.valid, 4) && ($past(in13.to, 4) == 15) && ($past(in13.data, 4) == out15.data) && (out15.from == 13)) || ($past(in14.valid, 4) && ($past(in14.to, 4) == 15) && ($past(in14.data, 4) == out15.data) && (out15.from == 14)) || ($past(in15.valid, 4) && ($past(in15.to, 4) == 15) && ($past(in15.data, 4) == out15.data) && (out15.from == 15)))));
    correct_output_exists: assert ((!$past(in0.valid, 4) || ((out0.valid && (out0.from == 0) && (out0.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 0)) || (out1.valid && (out1.from == 0) && (out1.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 1)) || (out2.valid && (out2.from == 0) && (out2.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 2)) || (out3.valid && (out3.from == 0) && (out3.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 3)) || (out4.valid && (out4.from == 0) && (out4.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 4)) || (out5.valid && (out5.from == 0) && (out5.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 5)) || (out6.valid && (out6.from == 0) && (out6.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 6)) || (out7.valid && (out7.from == 0) && (out7.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 7)) || (out8.valid && (out8.from == 0) && (out8.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 8)) || (out9.valid && (out9.from == 0) && (out9.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 9)) || (out10.valid && (out10.from == 0) && (out10.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 10)) || (out11.valid && (out11.from == 0) && (out11.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 11)) || (out12.valid && (out12.from == 0) && (out12.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 12)) || (out13.valid && (out13.from == 0) && (out13.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 13)) || (out14.valid && (out14.from == 0) && (out14.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 14)) || (out15.valid && (out15.from == 0) && (out15.data == $past(in0.data, 4)) && ($past(in0.to, 4) == 15))))
        && (!$past(in1.valid, 4) || ((out0.valid && (out0.from == 1) && (out0.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 0)) || (out1.valid && (out1.from == 1) && (out1.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 1)) || (out2.valid && (out2.from == 1) && (out2.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 2)) || (out3.valid && (out3.from == 1) && (out3.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 3)) || (out4.valid && (out4.from == 1) && (out4.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 4)) || (out5.valid && (out5.from == 1) && (out5.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 5)) || (out6.valid && (out6.from == 1) && (out6.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 6)) || (out7.valid && (out7.from == 1) && (out7.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 7)) || (out8.valid && (out8.from == 1) && (out8.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 8)) || (out9.valid && (out9.from == 1) && (out9.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 9)) || (out10.valid && (out10.from == 1) && (out10.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 10)) || (out11.valid && (out11.from == 1) && (out11.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 11)) || (out12.valid && (out12.from == 1) && (out12.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 12)) || (out13.valid && (out13.from == 1) && (out13.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 13)) || (out14.valid && (out14.from == 1) && (out14.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 14)) || (out15.valid && (out15.from == 1) && (out15.data == $past(in1.data, 4)) && ($past(in1.to, 4) == 15))))
        && (!$past(in2.valid, 4) || ((out0.valid && (out0.from == 2) && (out0.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 0)) || (out1.valid && (out1.from == 2) && (out1.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 1)) || (out2.valid && (out2.from == 2) && (out2.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 2)) || (out3.valid && (out3.from == 2) && (out3.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 3)) || (out4.valid && (out4.from == 2) && (out4.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 4)) || (out5.valid && (out5.from == 2) && (out5.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 5)) || (out6.valid && (out6.from == 2) && (out6.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 6)) || (out7.valid && (out7.from == 2) && (out7.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 7)) || (out8.valid && (out8.from == 2) && (out8.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 8)) || (out9.valid && (out9.from == 2) && (out9.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 9)) || (out10.valid && (out10.from == 2) && (out10.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 10)) || (out11.valid && (out11.from == 2) && (out11.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 11)) || (out12.valid && (out12.from == 2) && (out12.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 12)) || (out13.valid && (out13.from == 2) && (out13.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 13)) || (out14.valid && (out14.from == 2) && (out14.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 14)) || (out15.valid && (out15.from == 2) && (out15.data == $past(in2.data, 4)) && ($past(in2.to, 4) == 15))))
        && (!$past(in3.valid, 4) || ((out0.valid && (out0.from == 3) && (out0.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 0)) || (out1.valid && (out1.from == 3) && (out1.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 1)) || (out2.valid && (out2.from == 3) && (out2.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 2)) || (out3.valid && (out3.from == 3) && (out3.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 3)) || (out4.valid && (out4.from == 3) && (out4.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 4)) || (out5.valid && (out5.from == 3) && (out5.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 5)) || (out6.valid && (out6.from == 3) && (out6.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 6)) || (out7.valid && (out7.from == 3) && (out7.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 7)) || (out8.valid && (out8.from == 3) && (out8.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 8)) || (out9.valid && (out9.from == 3) && (out9.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 9)) || (out10.valid && (out10.from == 3) && (out10.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 10)) || (out11.valid && (out11.from == 3) && (out11.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 11)) || (out12.valid && (out12.from == 3) && (out12.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 12)) || (out13.valid && (out13.from == 3) && (out13.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 13)) || (out14.valid && (out14.from == 3) && (out14.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 14)) || (out15.valid && (out15.from == 3) && (out15.data == $past(in3.data, 4)) && ($past(in3.to, 4) == 15))))
        && (!$past(in4.valid, 4) || ((out0.valid && (out0.from == 4) && (out0.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 0)) || (out1.valid && (out1.from == 4) && (out1.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 1)) || (out2.valid && (out2.from == 4) && (out2.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 2)) || (out3.valid && (out3.from == 4) && (out3.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 3)) || (out4.valid && (out4.from == 4) && (out4.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 4)) || (out5.valid && (out5.from == 4) && (out5.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 5)) || (out6.valid && (out6.from == 4) && (out6.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 6)) || (out7.valid && (out7.from == 4) && (out7.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 7)) || (out8.valid && (out8.from == 4) && (out8.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 8)) || (out9.valid && (out9.from == 4) && (out9.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 9)) || (out10.valid && (out10.from == 4) && (out10.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 10)) || (out11.valid && (out11.from == 4) && (out11.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 11)) || (out12.valid && (out12.from == 4) && (out12.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 12)) || (out13.valid && (out13.from == 4) && (out13.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 13)) || (out14.valid && (out14.from == 4) && (out14.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 14)) || (out15.valid && (out15.from == 4) && (out15.data == $past(in4.data, 4)) && ($past(in4.to, 4) == 15))))
        && (!$past(in5.valid, 4) || ((out0.valid && (out0.from == 5) && (out0.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 0)) || (out1.valid && (out1.from == 5) && (out1.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 1)) || (out2.valid && (out2.from == 5) && (out2.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 2)) || (out3.valid && (out3.from == 5) && (out3.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 3)) || (out4.valid && (out4.from == 5) && (out4.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 4)) || (out5.valid && (out5.from == 5) && (out5.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 5)) || (out6.valid && (out6.from == 5) && (out6.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 6)) || (out7.valid && (out7.from == 5) && (out7.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 7)) || (out8.valid && (out8.from == 5) && (out8.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 8)) || (out9.valid && (out9.from == 5) && (out9.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 9)) || (out10.valid && (out10.from == 5) && (out10.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 10)) || (out11.valid && (out11.from == 5) && (out11.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 11)) || (out12.valid && (out12.from == 5) && (out12.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 12)) || (out13.valid && (out13.from == 5) && (out13.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 13)) || (out14.valid && (out14.from == 5) && (out14.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 14)) || (out15.valid && (out15.from == 5) && (out15.data == $past(in5.data, 4)) && ($past(in5.to, 4) == 15))))
        && (!$past(in6.valid, 4) || ((out0.valid && (out0.from == 6) && (out0.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 0)) || (out1.valid && (out1.from == 6) && (out1.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 1)) || (out2.valid && (out2.from == 6) && (out2.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 2)) || (out3.valid && (out3.from == 6) && (out3.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 3)) || (out4.valid && (out4.from == 6) && (out4.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 4)) || (out5.valid && (out5.from == 6) && (out5.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 5)) || (out6.valid && (out6.from == 6) && (out6.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 6)) || (out7.valid && (out7.from == 6) && (out7.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 7)) || (out8.valid && (out8.from == 6) && (out8.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 8)) || (out9.valid && (out9.from == 6) && (out9.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 9)) || (out10.valid && (out10.from == 6) && (out10.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 10)) || (out11.valid && (out11.from == 6) && (out11.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 11)) || (out12.valid && (out12.from == 6) && (out12.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 12)) || (out13.valid && (out13.from == 6) && (out13.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 13)) || (out14.valid && (out14.from == 6) && (out14.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 14)) || (out15.valid && (out15.from == 6) && (out15.data == $past(in6.data, 4)) && ($past(in6.to, 4) == 15))))
        && (!$past(in7.valid, 4) || ((out0.valid && (out0.from == 7) && (out0.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 0)) || (out1.valid && (out1.from == 7) && (out1.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 1)) || (out2.valid && (out2.from == 7) && (out2.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 2)) || (out3.valid && (out3.from == 7) && (out3.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 3)) || (out4.valid && (out4.from == 7) && (out4.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 4)) || (out5.valid && (out5.from == 7) && (out5.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 5)) || (out6.valid && (out6.from == 7) && (out6.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 6)) || (out7.valid && (out7.from == 7) && (out7.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 7)) || (out8.valid && (out8.from == 7) && (out8.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 8)) || (out9.valid && (out9.from == 7) && (out9.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 9)) || (out10.valid && (out10.from == 7) && (out10.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 10)) || (out11.valid && (out11.from == 7) && (out11.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 11)) || (out12.valid && (out12.from == 7) && (out12.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 12)) || (out13.valid && (out13.from == 7) && (out13.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 13)) || (out14.valid && (out14.from == 7) && (out14.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 14)) || (out15.valid && (out15.from == 7) && (out15.data == $past(in7.data, 4)) && ($past(in7.to, 4) == 15))))
        && (!$past(in8.valid, 4) || ((out0.valid && (out0.from == 8) && (out0.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 0)) || (out1.valid && (out1.from == 8) && (out1.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 1)) || (out2.valid && (out2.from == 8) && (out2.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 2)) || (out3.valid && (out3.from == 8) && (out3.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 3)) || (out4.valid && (out4.from == 8) && (out4.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 4)) || (out5.valid && (out5.from == 8) && (out5.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 5)) || (out6.valid && (out6.from == 8) && (out6.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 6)) || (out7.valid && (out7.from == 8) && (out7.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 7)) || (out8.valid && (out8.from == 8) && (out8.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 8)) || (out9.valid && (out9.from == 8) && (out9.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 9)) || (out10.valid && (out10.from == 8) && (out10.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 10)) || (out11.valid && (out11.from == 8) && (out11.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 11)) || (out12.valid && (out12.from == 8) && (out12.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 12)) || (out13.valid && (out13.from == 8) && (out13.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 13)) || (out14.valid && (out14.from == 8) && (out14.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 14)) || (out15.valid && (out15.from == 8) && (out15.data == $past(in8.data, 4)) && ($past(in8.to, 4) == 15))))
        && (!$past(in9.valid, 4) || ((out0.valid && (out0.from == 9) && (out0.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 0)) || (out1.valid && (out1.from == 9) && (out1.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 1)) || (out2.valid && (out2.from == 9) && (out2.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 2)) || (out3.valid && (out3.from == 9) && (out3.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 3)) || (out4.valid && (out4.from == 9) && (out4.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 4)) || (out5.valid && (out5.from == 9) && (out5.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 5)) || (out6.valid && (out6.from == 9) && (out6.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 6)) || (out7.valid && (out7.from == 9) && (out7.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 7)) || (out8.valid && (out8.from == 9) && (out8.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 8)) || (out9.valid && (out9.from == 9) && (out9.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 9)) || (out10.valid && (out10.from == 9) && (out10.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 10)) || (out11.valid && (out11.from == 9) && (out11.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 11)) || (out12.valid && (out12.from == 9) && (out12.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 12)) || (out13.valid && (out13.from == 9) && (out13.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 13)) || (out14.valid && (out14.from == 9) && (out14.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 14)) || (out15.valid && (out15.from == 9) && (out15.data == $past(in9.data, 4)) && ($past(in9.to, 4) == 15))))
        && (!$past(in10.valid, 4) || ((out0.valid && (out0.from == 10) && (out0.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 0)) || (out1.valid && (out1.from == 10) && (out1.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 1)) || (out2.valid && (out2.from == 10) && (out2.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 2)) || (out3.valid && (out3.from == 10) && (out3.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 3)) || (out4.valid && (out4.from == 10) && (out4.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 4)) || (out5.valid && (out5.from == 10) && (out5.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 5)) || (out6.valid && (out6.from == 10) && (out6.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 6)) || (out7.valid && (out7.from == 10) && (out7.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 7)) || (out8.valid && (out8.from == 10) && (out8.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 8)) || (out9.valid && (out9.from == 10) && (out9.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 9)) || (out10.valid && (out10.from == 10) && (out10.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 10)) || (out11.valid && (out11.from == 10) && (out11.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 11)) || (out12.valid && (out12.from == 10) && (out12.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 12)) || (out13.valid && (out13.from == 10) && (out13.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 13)) || (out14.valid && (out14.from == 10) && (out14.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 14)) || (out15.valid && (out15.from == 10) && (out15.data == $past(in10.data, 4)) && ($past(in10.to, 4) == 15))))
        && (!$past(in11.valid, 4) || ((out0.valid && (out0.from == 11) && (out0.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 0)) || (out1.valid && (out1.from == 11) && (out1.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 1)) || (out2.valid && (out2.from == 11) && (out2.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 2)) || (out3.valid && (out3.from == 11) && (out3.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 3)) || (out4.valid && (out4.from == 11) && (out4.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 4)) || (out5.valid && (out5.from == 11) && (out5.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 5)) || (out6.valid && (out6.from == 11) && (out6.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 6)) || (out7.valid && (out7.from == 11) && (out7.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 7)) || (out8.valid && (out8.from == 11) && (out8.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 8)) || (out9.valid && (out9.from == 11) && (out9.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 9)) || (out10.valid && (out10.from == 11) && (out10.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 10)) || (out11.valid && (out11.from == 11) && (out11.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 11)) || (out12.valid && (out12.from == 11) && (out12.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 12)) || (out13.valid && (out13.from == 11) && (out13.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 13)) || (out14.valid && (out14.from == 11) && (out14.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 14)) || (out15.valid && (out15.from == 11) && (out15.data == $past(in11.data, 4)) && ($past(in11.to, 4) == 15))))
        && (!$past(in12.valid, 4) || ((out0.valid && (out0.from == 12) && (out0.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 0)) || (out1.valid && (out1.from == 12) && (out1.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 1)) || (out2.valid && (out2.from == 12) && (out2.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 2)) || (out3.valid && (out3.from == 12) && (out3.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 3)) || (out4.valid && (out4.from == 12) && (out4.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 4)) || (out5.valid && (out5.from == 12) && (out5.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 5)) || (out6.valid && (out6.from == 12) && (out6.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 6)) || (out7.valid && (out7.from == 12) && (out7.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 7)) || (out8.valid && (out8.from == 12) && (out8.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 8)) || (out9.valid && (out9.from == 12) && (out9.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 9)) || (out10.valid && (out10.from == 12) && (out10.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 10)) || (out11.valid && (out11.from == 12) && (out11.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 11)) || (out12.valid && (out12.from == 12) && (out12.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 12)) || (out13.valid && (out13.from == 12) && (out13.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 13)) || (out14.valid && (out14.from == 12) && (out14.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 14)) || (out15.valid && (out15.from == 12) && (out15.data == $past(in12.data, 4)) && ($past(in12.to, 4) == 15))))
        && (!$past(in13.valid, 4) || ((out0.valid && (out0.from == 13) && (out0.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 0)) || (out1.valid && (out1.from == 13) && (out1.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 1)) || (out2.valid && (out2.from == 13) && (out2.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 2)) || (out3.valid && (out3.from == 13) && (out3.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 3)) || (out4.valid && (out4.from == 13) && (out4.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 4)) || (out5.valid && (out5.from == 13) && (out5.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 5)) || (out6.valid && (out6.from == 13) && (out6.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 6)) || (out7.valid && (out7.from == 13) && (out7.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 7)) || (out8.valid && (out8.from == 13) && (out8.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 8)) || (out9.valid && (out9.from == 13) && (out9.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 9)) || (out10.valid && (out10.from == 13) && (out10.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 10)) || (out11.valid && (out11.from == 13) && (out11.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 11)) || (out12.valid && (out12.from == 13) && (out12.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 12)) || (out13.valid && (out13.from == 13) && (out13.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 13)) || (out14.valid && (out14.from == 13) && (out14.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 14)) || (out15.valid && (out15.from == 13) && (out15.data == $past(in13.data, 4)) && ($past(in13.to, 4) == 15))))
        && (!$past(in14.valid, 4) || ((out0.valid && (out0.from == 14) && (out0.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 0)) || (out1.valid && (out1.from == 14) && (out1.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 1)) || (out2.valid && (out2.from == 14) && (out2.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 2)) || (out3.valid && (out3.from == 14) && (out3.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 3)) || (out4.valid && (out4.from == 14) && (out4.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 4)) || (out5.valid && (out5.from == 14) && (out5.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 5)) || (out6.valid && (out6.from == 14) && (out6.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 6)) || (out7.valid && (out7.from == 14) && (out7.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 7)) || (out8.valid && (out8.from == 14) && (out8.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 8)) || (out9.valid && (out9.from == 14) && (out9.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 9)) || (out10.valid && (out10.from == 14) && (out10.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 10)) || (out11.valid && (out11.from == 14) && (out11.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 11)) || (out12.valid && (out12.from == 14) && (out12.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 12)) || (out13.valid && (out13.from == 14) && (out13.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 13)) || (out14.valid && (out14.from == 14) && (out14.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 14)) || (out15.valid && (out15.from == 14) && (out15.data == $past(in14.data, 4)) && ($past(in14.to, 4) == 15))))
        && (!$past(in15.valid, 4) || ((out0.valid && (out0.from == 15) && (out0.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 0)) || (out1.valid && (out1.from == 15) && (out1.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 1)) || (out2.valid && (out2.from == 15) && (out2.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 2)) || (out3.valid && (out3.from == 15) && (out3.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 3)) || (out4.valid && (out4.from == 15) && (out4.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 4)) || (out5.valid && (out5.from == 15) && (out5.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 5)) || (out6.valid && (out6.from == 15) && (out6.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 6)) || (out7.valid && (out7.from == 15) && (out7.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 7)) || (out8.valid && (out8.from == 15) && (out8.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 8)) || (out9.valid && (out9.from == 15) && (out9.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 9)) || (out10.valid && (out10.from == 15) && (out10.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 10)) || (out11.valid && (out11.from == 15) && (out11.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 11)) || (out12.valid && (out12.from == 15) && (out12.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 12)) || (out13.valid && (out13.from == 15) && (out13.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 13)) || (out14.valid && (out14.from == 15) && (out14.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 14)) || (out15.valid && (out15.from == 15) && (out15.data == $past(in15.data, 4)) && ($past(in15.to, 4) == 15)))));
  end
end
`endif
endmodule
