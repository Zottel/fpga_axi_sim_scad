`default_nettype none

module TNT_BIN_HC0_JaSJ17_68_16_0 (
output wire [73-1:0] out0,
output wire [73-1:0] out1,
output wire [73-1:0] out2,
output wire [73-1:0] out3,
output wire [73-1:0] out4,
output wire [73-1:0] out5,
output wire [73-1:0] out6,
output wire [73-1:0] out7,
output wire [73-1:0] out8,
output wire [73-1:0] out9,
output wire [73-1:0] out10,
output wire [73-1:0] out11,
output wire [73-1:0] out12,
output wire [73-1:0] out13,
output wire [73-1:0] out14,
output wire [73-1:0] out15,
input wire [73-1:0] in0,
input wire [73-1:0] in1,
input wire [73-1:0] in2,
input wire [73-1:0] in3,
input wire [73-1:0] in4,
input wire [73-1:0] in5,
input wire [73-1:0] in6,
input wire [73-1:0] in7,
input wire [73-1:0] in8,
input wire [73-1:0] in9,
input wire [73-1:0] in10,
input wire [73-1:0] in11,
input wire [73-1:0] in12,
input wire [73-1:0] in13,
input wire [73-1:0] in14,
input wire [73-1:0] in15);
    wire x0_0;
    wire x0_1;
    wire x0_2;
    wire x0_3;
    wire x0_4;
    wire x0_5;
    wire x0_6;
    wire x0_7;
    wire x0_8;
    wire x0_9;
    wire x0_10;
    wire x0_11;
    wire x0_12;
    wire x0_13;
    wire x0_14;
    wire x0_15;
    wire x0_16;
    wire x0_17;
    wire x0_18;
    wire x0_19;
    wire x0_20;
    wire x0_21;
    wire x0_22;
    wire x0_23;
    wire x0_24;
    wire x0_25;
    wire x0_26;
    wire x0_27;
    wire x0_28;
    wire x0_29;
    wire x0_30;
    wire x0_31;
    wire x0_32;
    wire x0_33;
    wire x0_34;
    wire x0_35;
    wire x0_36;
    wire x0_37;
    wire x0_38;
    wire x0_39;
    wire x0_40;
    wire x0_41;
    wire x0_42;
    wire x0_43;
    wire x0_44;
    wire x0_45;
    wire x0_46;
    wire x0_47;
    wire x0_48;
    wire x0_49;
    wire x0_50;
    wire x0_51;
    wire x0_52;
    wire x0_53;
    wire x0_54;
    wire x0_55;
    wire x0_56;
    wire x0_57;
    wire x0_58;
    wire x0_59;
    wire x0_60;
    wire x0_61;
    wire x0_62;
    wire x0_63;
    wire x0_64;
    wire x0_65;
    wire x0_66;
    wire x0_67;
    wire x0_68;
    wire x0_69;
    wire x0_70;
    wire x0_71;
    wire x0_72;
    assign x0_0 = in0[0];
    assign x0_1 = in0[1];
    assign x0_2 = in0[2];
    assign x0_3 = in0[3];
    assign x0_4 = in0[4];
    assign x0_5 = in0[5];
    assign x0_6 = in0[6];
    assign x0_7 = in0[7];
    assign x0_8 = in0[8];
    assign x0_9 = in0[9];
    assign x0_10 = in0[10];
    assign x0_11 = in0[11];
    assign x0_12 = in0[12];
    assign x0_13 = in0[13];
    assign x0_14 = in0[14];
    assign x0_15 = in0[15];
    assign x0_16 = in0[16];
    assign x0_17 = in0[17];
    assign x0_18 = in0[18];
    assign x0_19 = in0[19];
    assign x0_20 = in0[20];
    assign x0_21 = in0[21];
    assign x0_22 = in0[22];
    assign x0_23 = in0[23];
    assign x0_24 = in0[24];
    assign x0_25 = in0[25];
    assign x0_26 = in0[26];
    assign x0_27 = in0[27];
    assign x0_28 = in0[28];
    assign x0_29 = in0[29];
    assign x0_30 = in0[30];
    assign x0_31 = in0[31];
    assign x0_32 = in0[32];
    assign x0_33 = in0[33];
    assign x0_34 = in0[34];
    assign x0_35 = in0[35];
    assign x0_36 = in0[36];
    assign x0_37 = in0[37];
    assign x0_38 = in0[38];
    assign x0_39 = in0[39];
    assign x0_40 = in0[40];
    assign x0_41 = in0[41];
    assign x0_42 = in0[42];
    assign x0_43 = in0[43];
    assign x0_44 = in0[44];
    assign x0_45 = in0[45];
    assign x0_46 = in0[46];
    assign x0_47 = in0[47];
    assign x0_48 = in0[48];
    assign x0_49 = in0[49];
    assign x0_50 = in0[50];
    assign x0_51 = in0[51];
    assign x0_52 = in0[52];
    assign x0_53 = in0[53];
    assign x0_54 = in0[54];
    assign x0_55 = in0[55];
    assign x0_56 = in0[56];
    assign x0_57 = in0[57];
    assign x0_58 = in0[58];
    assign x0_59 = in0[59];
    assign x0_60 = in0[60];
    assign x0_61 = in0[61];
    assign x0_62 = in0[62];
    assign x0_63 = in0[63];
    assign x0_64 = in0[64];
    assign x0_65 = in0[65];
    assign x0_66 = in0[66];
    assign x0_67 = in0[67];
    assign x0_68 = in0[68];
    assign x0_69 = in0[69];
    assign x0_70 = in0[70];
    assign x0_71 = in0[71];
    assign x0_72 = in0[72];
    wire x1_0;
    wire x1_1;
    wire x1_2;
    wire x1_3;
    wire x1_4;
    wire x1_5;
    wire x1_6;
    wire x1_7;
    wire x1_8;
    wire x1_9;
    wire x1_10;
    wire x1_11;
    wire x1_12;
    wire x1_13;
    wire x1_14;
    wire x1_15;
    wire x1_16;
    wire x1_17;
    wire x1_18;
    wire x1_19;
    wire x1_20;
    wire x1_21;
    wire x1_22;
    wire x1_23;
    wire x1_24;
    wire x1_25;
    wire x1_26;
    wire x1_27;
    wire x1_28;
    wire x1_29;
    wire x1_30;
    wire x1_31;
    wire x1_32;
    wire x1_33;
    wire x1_34;
    wire x1_35;
    wire x1_36;
    wire x1_37;
    wire x1_38;
    wire x1_39;
    wire x1_40;
    wire x1_41;
    wire x1_42;
    wire x1_43;
    wire x1_44;
    wire x1_45;
    wire x1_46;
    wire x1_47;
    wire x1_48;
    wire x1_49;
    wire x1_50;
    wire x1_51;
    wire x1_52;
    wire x1_53;
    wire x1_54;
    wire x1_55;
    wire x1_56;
    wire x1_57;
    wire x1_58;
    wire x1_59;
    wire x1_60;
    wire x1_61;
    wire x1_62;
    wire x1_63;
    wire x1_64;
    wire x1_65;
    wire x1_66;
    wire x1_67;
    wire x1_68;
    wire x1_69;
    wire x1_70;
    wire x1_71;
    wire x1_72;
    assign x1_0 = in1[0];
    assign x1_1 = in1[1];
    assign x1_2 = in1[2];
    assign x1_3 = in1[3];
    assign x1_4 = in1[4];
    assign x1_5 = in1[5];
    assign x1_6 = in1[6];
    assign x1_7 = in1[7];
    assign x1_8 = in1[8];
    assign x1_9 = in1[9];
    assign x1_10 = in1[10];
    assign x1_11 = in1[11];
    assign x1_12 = in1[12];
    assign x1_13 = in1[13];
    assign x1_14 = in1[14];
    assign x1_15 = in1[15];
    assign x1_16 = in1[16];
    assign x1_17 = in1[17];
    assign x1_18 = in1[18];
    assign x1_19 = in1[19];
    assign x1_20 = in1[20];
    assign x1_21 = in1[21];
    assign x1_22 = in1[22];
    assign x1_23 = in1[23];
    assign x1_24 = in1[24];
    assign x1_25 = in1[25];
    assign x1_26 = in1[26];
    assign x1_27 = in1[27];
    assign x1_28 = in1[28];
    assign x1_29 = in1[29];
    assign x1_30 = in1[30];
    assign x1_31 = in1[31];
    assign x1_32 = in1[32];
    assign x1_33 = in1[33];
    assign x1_34 = in1[34];
    assign x1_35 = in1[35];
    assign x1_36 = in1[36];
    assign x1_37 = in1[37];
    assign x1_38 = in1[38];
    assign x1_39 = in1[39];
    assign x1_40 = in1[40];
    assign x1_41 = in1[41];
    assign x1_42 = in1[42];
    assign x1_43 = in1[43];
    assign x1_44 = in1[44];
    assign x1_45 = in1[45];
    assign x1_46 = in1[46];
    assign x1_47 = in1[47];
    assign x1_48 = in1[48];
    assign x1_49 = in1[49];
    assign x1_50 = in1[50];
    assign x1_51 = in1[51];
    assign x1_52 = in1[52];
    assign x1_53 = in1[53];
    assign x1_54 = in1[54];
    assign x1_55 = in1[55];
    assign x1_56 = in1[56];
    assign x1_57 = in1[57];
    assign x1_58 = in1[58];
    assign x1_59 = in1[59];
    assign x1_60 = in1[60];
    assign x1_61 = in1[61];
    assign x1_62 = in1[62];
    assign x1_63 = in1[63];
    assign x1_64 = in1[64];
    assign x1_65 = in1[65];
    assign x1_66 = in1[66];
    assign x1_67 = in1[67];
    assign x1_68 = in1[68];
    assign x1_69 = in1[69];
    assign x1_70 = in1[70];
    assign x1_71 = in1[71];
    assign x1_72 = in1[72];
    wire x2_0;
    wire x2_1;
    wire x2_2;
    wire x2_3;
    wire x2_4;
    wire x2_5;
    wire x2_6;
    wire x2_7;
    wire x2_8;
    wire x2_9;
    wire x2_10;
    wire x2_11;
    wire x2_12;
    wire x2_13;
    wire x2_14;
    wire x2_15;
    wire x2_16;
    wire x2_17;
    wire x2_18;
    wire x2_19;
    wire x2_20;
    wire x2_21;
    wire x2_22;
    wire x2_23;
    wire x2_24;
    wire x2_25;
    wire x2_26;
    wire x2_27;
    wire x2_28;
    wire x2_29;
    wire x2_30;
    wire x2_31;
    wire x2_32;
    wire x2_33;
    wire x2_34;
    wire x2_35;
    wire x2_36;
    wire x2_37;
    wire x2_38;
    wire x2_39;
    wire x2_40;
    wire x2_41;
    wire x2_42;
    wire x2_43;
    wire x2_44;
    wire x2_45;
    wire x2_46;
    wire x2_47;
    wire x2_48;
    wire x2_49;
    wire x2_50;
    wire x2_51;
    wire x2_52;
    wire x2_53;
    wire x2_54;
    wire x2_55;
    wire x2_56;
    wire x2_57;
    wire x2_58;
    wire x2_59;
    wire x2_60;
    wire x2_61;
    wire x2_62;
    wire x2_63;
    wire x2_64;
    wire x2_65;
    wire x2_66;
    wire x2_67;
    wire x2_68;
    wire x2_69;
    wire x2_70;
    wire x2_71;
    wire x2_72;
    assign x2_0 = in2[0];
    assign x2_1 = in2[1];
    assign x2_2 = in2[2];
    assign x2_3 = in2[3];
    assign x2_4 = in2[4];
    assign x2_5 = in2[5];
    assign x2_6 = in2[6];
    assign x2_7 = in2[7];
    assign x2_8 = in2[8];
    assign x2_9 = in2[9];
    assign x2_10 = in2[10];
    assign x2_11 = in2[11];
    assign x2_12 = in2[12];
    assign x2_13 = in2[13];
    assign x2_14 = in2[14];
    assign x2_15 = in2[15];
    assign x2_16 = in2[16];
    assign x2_17 = in2[17];
    assign x2_18 = in2[18];
    assign x2_19 = in2[19];
    assign x2_20 = in2[20];
    assign x2_21 = in2[21];
    assign x2_22 = in2[22];
    assign x2_23 = in2[23];
    assign x2_24 = in2[24];
    assign x2_25 = in2[25];
    assign x2_26 = in2[26];
    assign x2_27 = in2[27];
    assign x2_28 = in2[28];
    assign x2_29 = in2[29];
    assign x2_30 = in2[30];
    assign x2_31 = in2[31];
    assign x2_32 = in2[32];
    assign x2_33 = in2[33];
    assign x2_34 = in2[34];
    assign x2_35 = in2[35];
    assign x2_36 = in2[36];
    assign x2_37 = in2[37];
    assign x2_38 = in2[38];
    assign x2_39 = in2[39];
    assign x2_40 = in2[40];
    assign x2_41 = in2[41];
    assign x2_42 = in2[42];
    assign x2_43 = in2[43];
    assign x2_44 = in2[44];
    assign x2_45 = in2[45];
    assign x2_46 = in2[46];
    assign x2_47 = in2[47];
    assign x2_48 = in2[48];
    assign x2_49 = in2[49];
    assign x2_50 = in2[50];
    assign x2_51 = in2[51];
    assign x2_52 = in2[52];
    assign x2_53 = in2[53];
    assign x2_54 = in2[54];
    assign x2_55 = in2[55];
    assign x2_56 = in2[56];
    assign x2_57 = in2[57];
    assign x2_58 = in2[58];
    assign x2_59 = in2[59];
    assign x2_60 = in2[60];
    assign x2_61 = in2[61];
    assign x2_62 = in2[62];
    assign x2_63 = in2[63];
    assign x2_64 = in2[64];
    assign x2_65 = in2[65];
    assign x2_66 = in2[66];
    assign x2_67 = in2[67];
    assign x2_68 = in2[68];
    assign x2_69 = in2[69];
    assign x2_70 = in2[70];
    assign x2_71 = in2[71];
    assign x2_72 = in2[72];
    wire x3_0;
    wire x3_1;
    wire x3_2;
    wire x3_3;
    wire x3_4;
    wire x3_5;
    wire x3_6;
    wire x3_7;
    wire x3_8;
    wire x3_9;
    wire x3_10;
    wire x3_11;
    wire x3_12;
    wire x3_13;
    wire x3_14;
    wire x3_15;
    wire x3_16;
    wire x3_17;
    wire x3_18;
    wire x3_19;
    wire x3_20;
    wire x3_21;
    wire x3_22;
    wire x3_23;
    wire x3_24;
    wire x3_25;
    wire x3_26;
    wire x3_27;
    wire x3_28;
    wire x3_29;
    wire x3_30;
    wire x3_31;
    wire x3_32;
    wire x3_33;
    wire x3_34;
    wire x3_35;
    wire x3_36;
    wire x3_37;
    wire x3_38;
    wire x3_39;
    wire x3_40;
    wire x3_41;
    wire x3_42;
    wire x3_43;
    wire x3_44;
    wire x3_45;
    wire x3_46;
    wire x3_47;
    wire x3_48;
    wire x3_49;
    wire x3_50;
    wire x3_51;
    wire x3_52;
    wire x3_53;
    wire x3_54;
    wire x3_55;
    wire x3_56;
    wire x3_57;
    wire x3_58;
    wire x3_59;
    wire x3_60;
    wire x3_61;
    wire x3_62;
    wire x3_63;
    wire x3_64;
    wire x3_65;
    wire x3_66;
    wire x3_67;
    wire x3_68;
    wire x3_69;
    wire x3_70;
    wire x3_71;
    wire x3_72;
    assign x3_0 = in3[0];
    assign x3_1 = in3[1];
    assign x3_2 = in3[2];
    assign x3_3 = in3[3];
    assign x3_4 = in3[4];
    assign x3_5 = in3[5];
    assign x3_6 = in3[6];
    assign x3_7 = in3[7];
    assign x3_8 = in3[8];
    assign x3_9 = in3[9];
    assign x3_10 = in3[10];
    assign x3_11 = in3[11];
    assign x3_12 = in3[12];
    assign x3_13 = in3[13];
    assign x3_14 = in3[14];
    assign x3_15 = in3[15];
    assign x3_16 = in3[16];
    assign x3_17 = in3[17];
    assign x3_18 = in3[18];
    assign x3_19 = in3[19];
    assign x3_20 = in3[20];
    assign x3_21 = in3[21];
    assign x3_22 = in3[22];
    assign x3_23 = in3[23];
    assign x3_24 = in3[24];
    assign x3_25 = in3[25];
    assign x3_26 = in3[26];
    assign x3_27 = in3[27];
    assign x3_28 = in3[28];
    assign x3_29 = in3[29];
    assign x3_30 = in3[30];
    assign x3_31 = in3[31];
    assign x3_32 = in3[32];
    assign x3_33 = in3[33];
    assign x3_34 = in3[34];
    assign x3_35 = in3[35];
    assign x3_36 = in3[36];
    assign x3_37 = in3[37];
    assign x3_38 = in3[38];
    assign x3_39 = in3[39];
    assign x3_40 = in3[40];
    assign x3_41 = in3[41];
    assign x3_42 = in3[42];
    assign x3_43 = in3[43];
    assign x3_44 = in3[44];
    assign x3_45 = in3[45];
    assign x3_46 = in3[46];
    assign x3_47 = in3[47];
    assign x3_48 = in3[48];
    assign x3_49 = in3[49];
    assign x3_50 = in3[50];
    assign x3_51 = in3[51];
    assign x3_52 = in3[52];
    assign x3_53 = in3[53];
    assign x3_54 = in3[54];
    assign x3_55 = in3[55];
    assign x3_56 = in3[56];
    assign x3_57 = in3[57];
    assign x3_58 = in3[58];
    assign x3_59 = in3[59];
    assign x3_60 = in3[60];
    assign x3_61 = in3[61];
    assign x3_62 = in3[62];
    assign x3_63 = in3[63];
    assign x3_64 = in3[64];
    assign x3_65 = in3[65];
    assign x3_66 = in3[66];
    assign x3_67 = in3[67];
    assign x3_68 = in3[68];
    assign x3_69 = in3[69];
    assign x3_70 = in3[70];
    assign x3_71 = in3[71];
    assign x3_72 = in3[72];
    wire x4_0;
    wire x4_1;
    wire x4_2;
    wire x4_3;
    wire x4_4;
    wire x4_5;
    wire x4_6;
    wire x4_7;
    wire x4_8;
    wire x4_9;
    wire x4_10;
    wire x4_11;
    wire x4_12;
    wire x4_13;
    wire x4_14;
    wire x4_15;
    wire x4_16;
    wire x4_17;
    wire x4_18;
    wire x4_19;
    wire x4_20;
    wire x4_21;
    wire x4_22;
    wire x4_23;
    wire x4_24;
    wire x4_25;
    wire x4_26;
    wire x4_27;
    wire x4_28;
    wire x4_29;
    wire x4_30;
    wire x4_31;
    wire x4_32;
    wire x4_33;
    wire x4_34;
    wire x4_35;
    wire x4_36;
    wire x4_37;
    wire x4_38;
    wire x4_39;
    wire x4_40;
    wire x4_41;
    wire x4_42;
    wire x4_43;
    wire x4_44;
    wire x4_45;
    wire x4_46;
    wire x4_47;
    wire x4_48;
    wire x4_49;
    wire x4_50;
    wire x4_51;
    wire x4_52;
    wire x4_53;
    wire x4_54;
    wire x4_55;
    wire x4_56;
    wire x4_57;
    wire x4_58;
    wire x4_59;
    wire x4_60;
    wire x4_61;
    wire x4_62;
    wire x4_63;
    wire x4_64;
    wire x4_65;
    wire x4_66;
    wire x4_67;
    wire x4_68;
    wire x4_69;
    wire x4_70;
    wire x4_71;
    wire x4_72;
    assign x4_0 = in4[0];
    assign x4_1 = in4[1];
    assign x4_2 = in4[2];
    assign x4_3 = in4[3];
    assign x4_4 = in4[4];
    assign x4_5 = in4[5];
    assign x4_6 = in4[6];
    assign x4_7 = in4[7];
    assign x4_8 = in4[8];
    assign x4_9 = in4[9];
    assign x4_10 = in4[10];
    assign x4_11 = in4[11];
    assign x4_12 = in4[12];
    assign x4_13 = in4[13];
    assign x4_14 = in4[14];
    assign x4_15 = in4[15];
    assign x4_16 = in4[16];
    assign x4_17 = in4[17];
    assign x4_18 = in4[18];
    assign x4_19 = in4[19];
    assign x4_20 = in4[20];
    assign x4_21 = in4[21];
    assign x4_22 = in4[22];
    assign x4_23 = in4[23];
    assign x4_24 = in4[24];
    assign x4_25 = in4[25];
    assign x4_26 = in4[26];
    assign x4_27 = in4[27];
    assign x4_28 = in4[28];
    assign x4_29 = in4[29];
    assign x4_30 = in4[30];
    assign x4_31 = in4[31];
    assign x4_32 = in4[32];
    assign x4_33 = in4[33];
    assign x4_34 = in4[34];
    assign x4_35 = in4[35];
    assign x4_36 = in4[36];
    assign x4_37 = in4[37];
    assign x4_38 = in4[38];
    assign x4_39 = in4[39];
    assign x4_40 = in4[40];
    assign x4_41 = in4[41];
    assign x4_42 = in4[42];
    assign x4_43 = in4[43];
    assign x4_44 = in4[44];
    assign x4_45 = in4[45];
    assign x4_46 = in4[46];
    assign x4_47 = in4[47];
    assign x4_48 = in4[48];
    assign x4_49 = in4[49];
    assign x4_50 = in4[50];
    assign x4_51 = in4[51];
    assign x4_52 = in4[52];
    assign x4_53 = in4[53];
    assign x4_54 = in4[54];
    assign x4_55 = in4[55];
    assign x4_56 = in4[56];
    assign x4_57 = in4[57];
    assign x4_58 = in4[58];
    assign x4_59 = in4[59];
    assign x4_60 = in4[60];
    assign x4_61 = in4[61];
    assign x4_62 = in4[62];
    assign x4_63 = in4[63];
    assign x4_64 = in4[64];
    assign x4_65 = in4[65];
    assign x4_66 = in4[66];
    assign x4_67 = in4[67];
    assign x4_68 = in4[68];
    assign x4_69 = in4[69];
    assign x4_70 = in4[70];
    assign x4_71 = in4[71];
    assign x4_72 = in4[72];
    wire x5_0;
    wire x5_1;
    wire x5_2;
    wire x5_3;
    wire x5_4;
    wire x5_5;
    wire x5_6;
    wire x5_7;
    wire x5_8;
    wire x5_9;
    wire x5_10;
    wire x5_11;
    wire x5_12;
    wire x5_13;
    wire x5_14;
    wire x5_15;
    wire x5_16;
    wire x5_17;
    wire x5_18;
    wire x5_19;
    wire x5_20;
    wire x5_21;
    wire x5_22;
    wire x5_23;
    wire x5_24;
    wire x5_25;
    wire x5_26;
    wire x5_27;
    wire x5_28;
    wire x5_29;
    wire x5_30;
    wire x5_31;
    wire x5_32;
    wire x5_33;
    wire x5_34;
    wire x5_35;
    wire x5_36;
    wire x5_37;
    wire x5_38;
    wire x5_39;
    wire x5_40;
    wire x5_41;
    wire x5_42;
    wire x5_43;
    wire x5_44;
    wire x5_45;
    wire x5_46;
    wire x5_47;
    wire x5_48;
    wire x5_49;
    wire x5_50;
    wire x5_51;
    wire x5_52;
    wire x5_53;
    wire x5_54;
    wire x5_55;
    wire x5_56;
    wire x5_57;
    wire x5_58;
    wire x5_59;
    wire x5_60;
    wire x5_61;
    wire x5_62;
    wire x5_63;
    wire x5_64;
    wire x5_65;
    wire x5_66;
    wire x5_67;
    wire x5_68;
    wire x5_69;
    wire x5_70;
    wire x5_71;
    wire x5_72;
    assign x5_0 = in5[0];
    assign x5_1 = in5[1];
    assign x5_2 = in5[2];
    assign x5_3 = in5[3];
    assign x5_4 = in5[4];
    assign x5_5 = in5[5];
    assign x5_6 = in5[6];
    assign x5_7 = in5[7];
    assign x5_8 = in5[8];
    assign x5_9 = in5[9];
    assign x5_10 = in5[10];
    assign x5_11 = in5[11];
    assign x5_12 = in5[12];
    assign x5_13 = in5[13];
    assign x5_14 = in5[14];
    assign x5_15 = in5[15];
    assign x5_16 = in5[16];
    assign x5_17 = in5[17];
    assign x5_18 = in5[18];
    assign x5_19 = in5[19];
    assign x5_20 = in5[20];
    assign x5_21 = in5[21];
    assign x5_22 = in5[22];
    assign x5_23 = in5[23];
    assign x5_24 = in5[24];
    assign x5_25 = in5[25];
    assign x5_26 = in5[26];
    assign x5_27 = in5[27];
    assign x5_28 = in5[28];
    assign x5_29 = in5[29];
    assign x5_30 = in5[30];
    assign x5_31 = in5[31];
    assign x5_32 = in5[32];
    assign x5_33 = in5[33];
    assign x5_34 = in5[34];
    assign x5_35 = in5[35];
    assign x5_36 = in5[36];
    assign x5_37 = in5[37];
    assign x5_38 = in5[38];
    assign x5_39 = in5[39];
    assign x5_40 = in5[40];
    assign x5_41 = in5[41];
    assign x5_42 = in5[42];
    assign x5_43 = in5[43];
    assign x5_44 = in5[44];
    assign x5_45 = in5[45];
    assign x5_46 = in5[46];
    assign x5_47 = in5[47];
    assign x5_48 = in5[48];
    assign x5_49 = in5[49];
    assign x5_50 = in5[50];
    assign x5_51 = in5[51];
    assign x5_52 = in5[52];
    assign x5_53 = in5[53];
    assign x5_54 = in5[54];
    assign x5_55 = in5[55];
    assign x5_56 = in5[56];
    assign x5_57 = in5[57];
    assign x5_58 = in5[58];
    assign x5_59 = in5[59];
    assign x5_60 = in5[60];
    assign x5_61 = in5[61];
    assign x5_62 = in5[62];
    assign x5_63 = in5[63];
    assign x5_64 = in5[64];
    assign x5_65 = in5[65];
    assign x5_66 = in5[66];
    assign x5_67 = in5[67];
    assign x5_68 = in5[68];
    assign x5_69 = in5[69];
    assign x5_70 = in5[70];
    assign x5_71 = in5[71];
    assign x5_72 = in5[72];
    wire x6_0;
    wire x6_1;
    wire x6_2;
    wire x6_3;
    wire x6_4;
    wire x6_5;
    wire x6_6;
    wire x6_7;
    wire x6_8;
    wire x6_9;
    wire x6_10;
    wire x6_11;
    wire x6_12;
    wire x6_13;
    wire x6_14;
    wire x6_15;
    wire x6_16;
    wire x6_17;
    wire x6_18;
    wire x6_19;
    wire x6_20;
    wire x6_21;
    wire x6_22;
    wire x6_23;
    wire x6_24;
    wire x6_25;
    wire x6_26;
    wire x6_27;
    wire x6_28;
    wire x6_29;
    wire x6_30;
    wire x6_31;
    wire x6_32;
    wire x6_33;
    wire x6_34;
    wire x6_35;
    wire x6_36;
    wire x6_37;
    wire x6_38;
    wire x6_39;
    wire x6_40;
    wire x6_41;
    wire x6_42;
    wire x6_43;
    wire x6_44;
    wire x6_45;
    wire x6_46;
    wire x6_47;
    wire x6_48;
    wire x6_49;
    wire x6_50;
    wire x6_51;
    wire x6_52;
    wire x6_53;
    wire x6_54;
    wire x6_55;
    wire x6_56;
    wire x6_57;
    wire x6_58;
    wire x6_59;
    wire x6_60;
    wire x6_61;
    wire x6_62;
    wire x6_63;
    wire x6_64;
    wire x6_65;
    wire x6_66;
    wire x6_67;
    wire x6_68;
    wire x6_69;
    wire x6_70;
    wire x6_71;
    wire x6_72;
    assign x6_0 = in6[0];
    assign x6_1 = in6[1];
    assign x6_2 = in6[2];
    assign x6_3 = in6[3];
    assign x6_4 = in6[4];
    assign x6_5 = in6[5];
    assign x6_6 = in6[6];
    assign x6_7 = in6[7];
    assign x6_8 = in6[8];
    assign x6_9 = in6[9];
    assign x6_10 = in6[10];
    assign x6_11 = in6[11];
    assign x6_12 = in6[12];
    assign x6_13 = in6[13];
    assign x6_14 = in6[14];
    assign x6_15 = in6[15];
    assign x6_16 = in6[16];
    assign x6_17 = in6[17];
    assign x6_18 = in6[18];
    assign x6_19 = in6[19];
    assign x6_20 = in6[20];
    assign x6_21 = in6[21];
    assign x6_22 = in6[22];
    assign x6_23 = in6[23];
    assign x6_24 = in6[24];
    assign x6_25 = in6[25];
    assign x6_26 = in6[26];
    assign x6_27 = in6[27];
    assign x6_28 = in6[28];
    assign x6_29 = in6[29];
    assign x6_30 = in6[30];
    assign x6_31 = in6[31];
    assign x6_32 = in6[32];
    assign x6_33 = in6[33];
    assign x6_34 = in6[34];
    assign x6_35 = in6[35];
    assign x6_36 = in6[36];
    assign x6_37 = in6[37];
    assign x6_38 = in6[38];
    assign x6_39 = in6[39];
    assign x6_40 = in6[40];
    assign x6_41 = in6[41];
    assign x6_42 = in6[42];
    assign x6_43 = in6[43];
    assign x6_44 = in6[44];
    assign x6_45 = in6[45];
    assign x6_46 = in6[46];
    assign x6_47 = in6[47];
    assign x6_48 = in6[48];
    assign x6_49 = in6[49];
    assign x6_50 = in6[50];
    assign x6_51 = in6[51];
    assign x6_52 = in6[52];
    assign x6_53 = in6[53];
    assign x6_54 = in6[54];
    assign x6_55 = in6[55];
    assign x6_56 = in6[56];
    assign x6_57 = in6[57];
    assign x6_58 = in6[58];
    assign x6_59 = in6[59];
    assign x6_60 = in6[60];
    assign x6_61 = in6[61];
    assign x6_62 = in6[62];
    assign x6_63 = in6[63];
    assign x6_64 = in6[64];
    assign x6_65 = in6[65];
    assign x6_66 = in6[66];
    assign x6_67 = in6[67];
    assign x6_68 = in6[68];
    assign x6_69 = in6[69];
    assign x6_70 = in6[70];
    assign x6_71 = in6[71];
    assign x6_72 = in6[72];
    wire x7_0;
    wire x7_1;
    wire x7_2;
    wire x7_3;
    wire x7_4;
    wire x7_5;
    wire x7_6;
    wire x7_7;
    wire x7_8;
    wire x7_9;
    wire x7_10;
    wire x7_11;
    wire x7_12;
    wire x7_13;
    wire x7_14;
    wire x7_15;
    wire x7_16;
    wire x7_17;
    wire x7_18;
    wire x7_19;
    wire x7_20;
    wire x7_21;
    wire x7_22;
    wire x7_23;
    wire x7_24;
    wire x7_25;
    wire x7_26;
    wire x7_27;
    wire x7_28;
    wire x7_29;
    wire x7_30;
    wire x7_31;
    wire x7_32;
    wire x7_33;
    wire x7_34;
    wire x7_35;
    wire x7_36;
    wire x7_37;
    wire x7_38;
    wire x7_39;
    wire x7_40;
    wire x7_41;
    wire x7_42;
    wire x7_43;
    wire x7_44;
    wire x7_45;
    wire x7_46;
    wire x7_47;
    wire x7_48;
    wire x7_49;
    wire x7_50;
    wire x7_51;
    wire x7_52;
    wire x7_53;
    wire x7_54;
    wire x7_55;
    wire x7_56;
    wire x7_57;
    wire x7_58;
    wire x7_59;
    wire x7_60;
    wire x7_61;
    wire x7_62;
    wire x7_63;
    wire x7_64;
    wire x7_65;
    wire x7_66;
    wire x7_67;
    wire x7_68;
    wire x7_69;
    wire x7_70;
    wire x7_71;
    wire x7_72;
    assign x7_0 = in7[0];
    assign x7_1 = in7[1];
    assign x7_2 = in7[2];
    assign x7_3 = in7[3];
    assign x7_4 = in7[4];
    assign x7_5 = in7[5];
    assign x7_6 = in7[6];
    assign x7_7 = in7[7];
    assign x7_8 = in7[8];
    assign x7_9 = in7[9];
    assign x7_10 = in7[10];
    assign x7_11 = in7[11];
    assign x7_12 = in7[12];
    assign x7_13 = in7[13];
    assign x7_14 = in7[14];
    assign x7_15 = in7[15];
    assign x7_16 = in7[16];
    assign x7_17 = in7[17];
    assign x7_18 = in7[18];
    assign x7_19 = in7[19];
    assign x7_20 = in7[20];
    assign x7_21 = in7[21];
    assign x7_22 = in7[22];
    assign x7_23 = in7[23];
    assign x7_24 = in7[24];
    assign x7_25 = in7[25];
    assign x7_26 = in7[26];
    assign x7_27 = in7[27];
    assign x7_28 = in7[28];
    assign x7_29 = in7[29];
    assign x7_30 = in7[30];
    assign x7_31 = in7[31];
    assign x7_32 = in7[32];
    assign x7_33 = in7[33];
    assign x7_34 = in7[34];
    assign x7_35 = in7[35];
    assign x7_36 = in7[36];
    assign x7_37 = in7[37];
    assign x7_38 = in7[38];
    assign x7_39 = in7[39];
    assign x7_40 = in7[40];
    assign x7_41 = in7[41];
    assign x7_42 = in7[42];
    assign x7_43 = in7[43];
    assign x7_44 = in7[44];
    assign x7_45 = in7[45];
    assign x7_46 = in7[46];
    assign x7_47 = in7[47];
    assign x7_48 = in7[48];
    assign x7_49 = in7[49];
    assign x7_50 = in7[50];
    assign x7_51 = in7[51];
    assign x7_52 = in7[52];
    assign x7_53 = in7[53];
    assign x7_54 = in7[54];
    assign x7_55 = in7[55];
    assign x7_56 = in7[56];
    assign x7_57 = in7[57];
    assign x7_58 = in7[58];
    assign x7_59 = in7[59];
    assign x7_60 = in7[60];
    assign x7_61 = in7[61];
    assign x7_62 = in7[62];
    assign x7_63 = in7[63];
    assign x7_64 = in7[64];
    assign x7_65 = in7[65];
    assign x7_66 = in7[66];
    assign x7_67 = in7[67];
    assign x7_68 = in7[68];
    assign x7_69 = in7[69];
    assign x7_70 = in7[70];
    assign x7_71 = in7[71];
    assign x7_72 = in7[72];
    wire x8_0;
    wire x8_1;
    wire x8_2;
    wire x8_3;
    wire x8_4;
    wire x8_5;
    wire x8_6;
    wire x8_7;
    wire x8_8;
    wire x8_9;
    wire x8_10;
    wire x8_11;
    wire x8_12;
    wire x8_13;
    wire x8_14;
    wire x8_15;
    wire x8_16;
    wire x8_17;
    wire x8_18;
    wire x8_19;
    wire x8_20;
    wire x8_21;
    wire x8_22;
    wire x8_23;
    wire x8_24;
    wire x8_25;
    wire x8_26;
    wire x8_27;
    wire x8_28;
    wire x8_29;
    wire x8_30;
    wire x8_31;
    wire x8_32;
    wire x8_33;
    wire x8_34;
    wire x8_35;
    wire x8_36;
    wire x8_37;
    wire x8_38;
    wire x8_39;
    wire x8_40;
    wire x8_41;
    wire x8_42;
    wire x8_43;
    wire x8_44;
    wire x8_45;
    wire x8_46;
    wire x8_47;
    wire x8_48;
    wire x8_49;
    wire x8_50;
    wire x8_51;
    wire x8_52;
    wire x8_53;
    wire x8_54;
    wire x8_55;
    wire x8_56;
    wire x8_57;
    wire x8_58;
    wire x8_59;
    wire x8_60;
    wire x8_61;
    wire x8_62;
    wire x8_63;
    wire x8_64;
    wire x8_65;
    wire x8_66;
    wire x8_67;
    wire x8_68;
    wire x8_69;
    wire x8_70;
    wire x8_71;
    wire x8_72;
    assign x8_0 = in8[0];
    assign x8_1 = in8[1];
    assign x8_2 = in8[2];
    assign x8_3 = in8[3];
    assign x8_4 = in8[4];
    assign x8_5 = in8[5];
    assign x8_6 = in8[6];
    assign x8_7 = in8[7];
    assign x8_8 = in8[8];
    assign x8_9 = in8[9];
    assign x8_10 = in8[10];
    assign x8_11 = in8[11];
    assign x8_12 = in8[12];
    assign x8_13 = in8[13];
    assign x8_14 = in8[14];
    assign x8_15 = in8[15];
    assign x8_16 = in8[16];
    assign x8_17 = in8[17];
    assign x8_18 = in8[18];
    assign x8_19 = in8[19];
    assign x8_20 = in8[20];
    assign x8_21 = in8[21];
    assign x8_22 = in8[22];
    assign x8_23 = in8[23];
    assign x8_24 = in8[24];
    assign x8_25 = in8[25];
    assign x8_26 = in8[26];
    assign x8_27 = in8[27];
    assign x8_28 = in8[28];
    assign x8_29 = in8[29];
    assign x8_30 = in8[30];
    assign x8_31 = in8[31];
    assign x8_32 = in8[32];
    assign x8_33 = in8[33];
    assign x8_34 = in8[34];
    assign x8_35 = in8[35];
    assign x8_36 = in8[36];
    assign x8_37 = in8[37];
    assign x8_38 = in8[38];
    assign x8_39 = in8[39];
    assign x8_40 = in8[40];
    assign x8_41 = in8[41];
    assign x8_42 = in8[42];
    assign x8_43 = in8[43];
    assign x8_44 = in8[44];
    assign x8_45 = in8[45];
    assign x8_46 = in8[46];
    assign x8_47 = in8[47];
    assign x8_48 = in8[48];
    assign x8_49 = in8[49];
    assign x8_50 = in8[50];
    assign x8_51 = in8[51];
    assign x8_52 = in8[52];
    assign x8_53 = in8[53];
    assign x8_54 = in8[54];
    assign x8_55 = in8[55];
    assign x8_56 = in8[56];
    assign x8_57 = in8[57];
    assign x8_58 = in8[58];
    assign x8_59 = in8[59];
    assign x8_60 = in8[60];
    assign x8_61 = in8[61];
    assign x8_62 = in8[62];
    assign x8_63 = in8[63];
    assign x8_64 = in8[64];
    assign x8_65 = in8[65];
    assign x8_66 = in8[66];
    assign x8_67 = in8[67];
    assign x8_68 = in8[68];
    assign x8_69 = in8[69];
    assign x8_70 = in8[70];
    assign x8_71 = in8[71];
    assign x8_72 = in8[72];
    wire x9_0;
    wire x9_1;
    wire x9_2;
    wire x9_3;
    wire x9_4;
    wire x9_5;
    wire x9_6;
    wire x9_7;
    wire x9_8;
    wire x9_9;
    wire x9_10;
    wire x9_11;
    wire x9_12;
    wire x9_13;
    wire x9_14;
    wire x9_15;
    wire x9_16;
    wire x9_17;
    wire x9_18;
    wire x9_19;
    wire x9_20;
    wire x9_21;
    wire x9_22;
    wire x9_23;
    wire x9_24;
    wire x9_25;
    wire x9_26;
    wire x9_27;
    wire x9_28;
    wire x9_29;
    wire x9_30;
    wire x9_31;
    wire x9_32;
    wire x9_33;
    wire x9_34;
    wire x9_35;
    wire x9_36;
    wire x9_37;
    wire x9_38;
    wire x9_39;
    wire x9_40;
    wire x9_41;
    wire x9_42;
    wire x9_43;
    wire x9_44;
    wire x9_45;
    wire x9_46;
    wire x9_47;
    wire x9_48;
    wire x9_49;
    wire x9_50;
    wire x9_51;
    wire x9_52;
    wire x9_53;
    wire x9_54;
    wire x9_55;
    wire x9_56;
    wire x9_57;
    wire x9_58;
    wire x9_59;
    wire x9_60;
    wire x9_61;
    wire x9_62;
    wire x9_63;
    wire x9_64;
    wire x9_65;
    wire x9_66;
    wire x9_67;
    wire x9_68;
    wire x9_69;
    wire x9_70;
    wire x9_71;
    wire x9_72;
    assign x9_0 = in9[0];
    assign x9_1 = in9[1];
    assign x9_2 = in9[2];
    assign x9_3 = in9[3];
    assign x9_4 = in9[4];
    assign x9_5 = in9[5];
    assign x9_6 = in9[6];
    assign x9_7 = in9[7];
    assign x9_8 = in9[8];
    assign x9_9 = in9[9];
    assign x9_10 = in9[10];
    assign x9_11 = in9[11];
    assign x9_12 = in9[12];
    assign x9_13 = in9[13];
    assign x9_14 = in9[14];
    assign x9_15 = in9[15];
    assign x9_16 = in9[16];
    assign x9_17 = in9[17];
    assign x9_18 = in9[18];
    assign x9_19 = in9[19];
    assign x9_20 = in9[20];
    assign x9_21 = in9[21];
    assign x9_22 = in9[22];
    assign x9_23 = in9[23];
    assign x9_24 = in9[24];
    assign x9_25 = in9[25];
    assign x9_26 = in9[26];
    assign x9_27 = in9[27];
    assign x9_28 = in9[28];
    assign x9_29 = in9[29];
    assign x9_30 = in9[30];
    assign x9_31 = in9[31];
    assign x9_32 = in9[32];
    assign x9_33 = in9[33];
    assign x9_34 = in9[34];
    assign x9_35 = in9[35];
    assign x9_36 = in9[36];
    assign x9_37 = in9[37];
    assign x9_38 = in9[38];
    assign x9_39 = in9[39];
    assign x9_40 = in9[40];
    assign x9_41 = in9[41];
    assign x9_42 = in9[42];
    assign x9_43 = in9[43];
    assign x9_44 = in9[44];
    assign x9_45 = in9[45];
    assign x9_46 = in9[46];
    assign x9_47 = in9[47];
    assign x9_48 = in9[48];
    assign x9_49 = in9[49];
    assign x9_50 = in9[50];
    assign x9_51 = in9[51];
    assign x9_52 = in9[52];
    assign x9_53 = in9[53];
    assign x9_54 = in9[54];
    assign x9_55 = in9[55];
    assign x9_56 = in9[56];
    assign x9_57 = in9[57];
    assign x9_58 = in9[58];
    assign x9_59 = in9[59];
    assign x9_60 = in9[60];
    assign x9_61 = in9[61];
    assign x9_62 = in9[62];
    assign x9_63 = in9[63];
    assign x9_64 = in9[64];
    assign x9_65 = in9[65];
    assign x9_66 = in9[66];
    assign x9_67 = in9[67];
    assign x9_68 = in9[68];
    assign x9_69 = in9[69];
    assign x9_70 = in9[70];
    assign x9_71 = in9[71];
    assign x9_72 = in9[72];
    wire x10_0;
    wire x10_1;
    wire x10_2;
    wire x10_3;
    wire x10_4;
    wire x10_5;
    wire x10_6;
    wire x10_7;
    wire x10_8;
    wire x10_9;
    wire x10_10;
    wire x10_11;
    wire x10_12;
    wire x10_13;
    wire x10_14;
    wire x10_15;
    wire x10_16;
    wire x10_17;
    wire x10_18;
    wire x10_19;
    wire x10_20;
    wire x10_21;
    wire x10_22;
    wire x10_23;
    wire x10_24;
    wire x10_25;
    wire x10_26;
    wire x10_27;
    wire x10_28;
    wire x10_29;
    wire x10_30;
    wire x10_31;
    wire x10_32;
    wire x10_33;
    wire x10_34;
    wire x10_35;
    wire x10_36;
    wire x10_37;
    wire x10_38;
    wire x10_39;
    wire x10_40;
    wire x10_41;
    wire x10_42;
    wire x10_43;
    wire x10_44;
    wire x10_45;
    wire x10_46;
    wire x10_47;
    wire x10_48;
    wire x10_49;
    wire x10_50;
    wire x10_51;
    wire x10_52;
    wire x10_53;
    wire x10_54;
    wire x10_55;
    wire x10_56;
    wire x10_57;
    wire x10_58;
    wire x10_59;
    wire x10_60;
    wire x10_61;
    wire x10_62;
    wire x10_63;
    wire x10_64;
    wire x10_65;
    wire x10_66;
    wire x10_67;
    wire x10_68;
    wire x10_69;
    wire x10_70;
    wire x10_71;
    wire x10_72;
    assign x10_0 = in10[0];
    assign x10_1 = in10[1];
    assign x10_2 = in10[2];
    assign x10_3 = in10[3];
    assign x10_4 = in10[4];
    assign x10_5 = in10[5];
    assign x10_6 = in10[6];
    assign x10_7 = in10[7];
    assign x10_8 = in10[8];
    assign x10_9 = in10[9];
    assign x10_10 = in10[10];
    assign x10_11 = in10[11];
    assign x10_12 = in10[12];
    assign x10_13 = in10[13];
    assign x10_14 = in10[14];
    assign x10_15 = in10[15];
    assign x10_16 = in10[16];
    assign x10_17 = in10[17];
    assign x10_18 = in10[18];
    assign x10_19 = in10[19];
    assign x10_20 = in10[20];
    assign x10_21 = in10[21];
    assign x10_22 = in10[22];
    assign x10_23 = in10[23];
    assign x10_24 = in10[24];
    assign x10_25 = in10[25];
    assign x10_26 = in10[26];
    assign x10_27 = in10[27];
    assign x10_28 = in10[28];
    assign x10_29 = in10[29];
    assign x10_30 = in10[30];
    assign x10_31 = in10[31];
    assign x10_32 = in10[32];
    assign x10_33 = in10[33];
    assign x10_34 = in10[34];
    assign x10_35 = in10[35];
    assign x10_36 = in10[36];
    assign x10_37 = in10[37];
    assign x10_38 = in10[38];
    assign x10_39 = in10[39];
    assign x10_40 = in10[40];
    assign x10_41 = in10[41];
    assign x10_42 = in10[42];
    assign x10_43 = in10[43];
    assign x10_44 = in10[44];
    assign x10_45 = in10[45];
    assign x10_46 = in10[46];
    assign x10_47 = in10[47];
    assign x10_48 = in10[48];
    assign x10_49 = in10[49];
    assign x10_50 = in10[50];
    assign x10_51 = in10[51];
    assign x10_52 = in10[52];
    assign x10_53 = in10[53];
    assign x10_54 = in10[54];
    assign x10_55 = in10[55];
    assign x10_56 = in10[56];
    assign x10_57 = in10[57];
    assign x10_58 = in10[58];
    assign x10_59 = in10[59];
    assign x10_60 = in10[60];
    assign x10_61 = in10[61];
    assign x10_62 = in10[62];
    assign x10_63 = in10[63];
    assign x10_64 = in10[64];
    assign x10_65 = in10[65];
    assign x10_66 = in10[66];
    assign x10_67 = in10[67];
    assign x10_68 = in10[68];
    assign x10_69 = in10[69];
    assign x10_70 = in10[70];
    assign x10_71 = in10[71];
    assign x10_72 = in10[72];
    wire x11_0;
    wire x11_1;
    wire x11_2;
    wire x11_3;
    wire x11_4;
    wire x11_5;
    wire x11_6;
    wire x11_7;
    wire x11_8;
    wire x11_9;
    wire x11_10;
    wire x11_11;
    wire x11_12;
    wire x11_13;
    wire x11_14;
    wire x11_15;
    wire x11_16;
    wire x11_17;
    wire x11_18;
    wire x11_19;
    wire x11_20;
    wire x11_21;
    wire x11_22;
    wire x11_23;
    wire x11_24;
    wire x11_25;
    wire x11_26;
    wire x11_27;
    wire x11_28;
    wire x11_29;
    wire x11_30;
    wire x11_31;
    wire x11_32;
    wire x11_33;
    wire x11_34;
    wire x11_35;
    wire x11_36;
    wire x11_37;
    wire x11_38;
    wire x11_39;
    wire x11_40;
    wire x11_41;
    wire x11_42;
    wire x11_43;
    wire x11_44;
    wire x11_45;
    wire x11_46;
    wire x11_47;
    wire x11_48;
    wire x11_49;
    wire x11_50;
    wire x11_51;
    wire x11_52;
    wire x11_53;
    wire x11_54;
    wire x11_55;
    wire x11_56;
    wire x11_57;
    wire x11_58;
    wire x11_59;
    wire x11_60;
    wire x11_61;
    wire x11_62;
    wire x11_63;
    wire x11_64;
    wire x11_65;
    wire x11_66;
    wire x11_67;
    wire x11_68;
    wire x11_69;
    wire x11_70;
    wire x11_71;
    wire x11_72;
    assign x11_0 = in11[0];
    assign x11_1 = in11[1];
    assign x11_2 = in11[2];
    assign x11_3 = in11[3];
    assign x11_4 = in11[4];
    assign x11_5 = in11[5];
    assign x11_6 = in11[6];
    assign x11_7 = in11[7];
    assign x11_8 = in11[8];
    assign x11_9 = in11[9];
    assign x11_10 = in11[10];
    assign x11_11 = in11[11];
    assign x11_12 = in11[12];
    assign x11_13 = in11[13];
    assign x11_14 = in11[14];
    assign x11_15 = in11[15];
    assign x11_16 = in11[16];
    assign x11_17 = in11[17];
    assign x11_18 = in11[18];
    assign x11_19 = in11[19];
    assign x11_20 = in11[20];
    assign x11_21 = in11[21];
    assign x11_22 = in11[22];
    assign x11_23 = in11[23];
    assign x11_24 = in11[24];
    assign x11_25 = in11[25];
    assign x11_26 = in11[26];
    assign x11_27 = in11[27];
    assign x11_28 = in11[28];
    assign x11_29 = in11[29];
    assign x11_30 = in11[30];
    assign x11_31 = in11[31];
    assign x11_32 = in11[32];
    assign x11_33 = in11[33];
    assign x11_34 = in11[34];
    assign x11_35 = in11[35];
    assign x11_36 = in11[36];
    assign x11_37 = in11[37];
    assign x11_38 = in11[38];
    assign x11_39 = in11[39];
    assign x11_40 = in11[40];
    assign x11_41 = in11[41];
    assign x11_42 = in11[42];
    assign x11_43 = in11[43];
    assign x11_44 = in11[44];
    assign x11_45 = in11[45];
    assign x11_46 = in11[46];
    assign x11_47 = in11[47];
    assign x11_48 = in11[48];
    assign x11_49 = in11[49];
    assign x11_50 = in11[50];
    assign x11_51 = in11[51];
    assign x11_52 = in11[52];
    assign x11_53 = in11[53];
    assign x11_54 = in11[54];
    assign x11_55 = in11[55];
    assign x11_56 = in11[56];
    assign x11_57 = in11[57];
    assign x11_58 = in11[58];
    assign x11_59 = in11[59];
    assign x11_60 = in11[60];
    assign x11_61 = in11[61];
    assign x11_62 = in11[62];
    assign x11_63 = in11[63];
    assign x11_64 = in11[64];
    assign x11_65 = in11[65];
    assign x11_66 = in11[66];
    assign x11_67 = in11[67];
    assign x11_68 = in11[68];
    assign x11_69 = in11[69];
    assign x11_70 = in11[70];
    assign x11_71 = in11[71];
    assign x11_72 = in11[72];
    wire x12_0;
    wire x12_1;
    wire x12_2;
    wire x12_3;
    wire x12_4;
    wire x12_5;
    wire x12_6;
    wire x12_7;
    wire x12_8;
    wire x12_9;
    wire x12_10;
    wire x12_11;
    wire x12_12;
    wire x12_13;
    wire x12_14;
    wire x12_15;
    wire x12_16;
    wire x12_17;
    wire x12_18;
    wire x12_19;
    wire x12_20;
    wire x12_21;
    wire x12_22;
    wire x12_23;
    wire x12_24;
    wire x12_25;
    wire x12_26;
    wire x12_27;
    wire x12_28;
    wire x12_29;
    wire x12_30;
    wire x12_31;
    wire x12_32;
    wire x12_33;
    wire x12_34;
    wire x12_35;
    wire x12_36;
    wire x12_37;
    wire x12_38;
    wire x12_39;
    wire x12_40;
    wire x12_41;
    wire x12_42;
    wire x12_43;
    wire x12_44;
    wire x12_45;
    wire x12_46;
    wire x12_47;
    wire x12_48;
    wire x12_49;
    wire x12_50;
    wire x12_51;
    wire x12_52;
    wire x12_53;
    wire x12_54;
    wire x12_55;
    wire x12_56;
    wire x12_57;
    wire x12_58;
    wire x12_59;
    wire x12_60;
    wire x12_61;
    wire x12_62;
    wire x12_63;
    wire x12_64;
    wire x12_65;
    wire x12_66;
    wire x12_67;
    wire x12_68;
    wire x12_69;
    wire x12_70;
    wire x12_71;
    wire x12_72;
    assign x12_0 = in12[0];
    assign x12_1 = in12[1];
    assign x12_2 = in12[2];
    assign x12_3 = in12[3];
    assign x12_4 = in12[4];
    assign x12_5 = in12[5];
    assign x12_6 = in12[6];
    assign x12_7 = in12[7];
    assign x12_8 = in12[8];
    assign x12_9 = in12[9];
    assign x12_10 = in12[10];
    assign x12_11 = in12[11];
    assign x12_12 = in12[12];
    assign x12_13 = in12[13];
    assign x12_14 = in12[14];
    assign x12_15 = in12[15];
    assign x12_16 = in12[16];
    assign x12_17 = in12[17];
    assign x12_18 = in12[18];
    assign x12_19 = in12[19];
    assign x12_20 = in12[20];
    assign x12_21 = in12[21];
    assign x12_22 = in12[22];
    assign x12_23 = in12[23];
    assign x12_24 = in12[24];
    assign x12_25 = in12[25];
    assign x12_26 = in12[26];
    assign x12_27 = in12[27];
    assign x12_28 = in12[28];
    assign x12_29 = in12[29];
    assign x12_30 = in12[30];
    assign x12_31 = in12[31];
    assign x12_32 = in12[32];
    assign x12_33 = in12[33];
    assign x12_34 = in12[34];
    assign x12_35 = in12[35];
    assign x12_36 = in12[36];
    assign x12_37 = in12[37];
    assign x12_38 = in12[38];
    assign x12_39 = in12[39];
    assign x12_40 = in12[40];
    assign x12_41 = in12[41];
    assign x12_42 = in12[42];
    assign x12_43 = in12[43];
    assign x12_44 = in12[44];
    assign x12_45 = in12[45];
    assign x12_46 = in12[46];
    assign x12_47 = in12[47];
    assign x12_48 = in12[48];
    assign x12_49 = in12[49];
    assign x12_50 = in12[50];
    assign x12_51 = in12[51];
    assign x12_52 = in12[52];
    assign x12_53 = in12[53];
    assign x12_54 = in12[54];
    assign x12_55 = in12[55];
    assign x12_56 = in12[56];
    assign x12_57 = in12[57];
    assign x12_58 = in12[58];
    assign x12_59 = in12[59];
    assign x12_60 = in12[60];
    assign x12_61 = in12[61];
    assign x12_62 = in12[62];
    assign x12_63 = in12[63];
    assign x12_64 = in12[64];
    assign x12_65 = in12[65];
    assign x12_66 = in12[66];
    assign x12_67 = in12[67];
    assign x12_68 = in12[68];
    assign x12_69 = in12[69];
    assign x12_70 = in12[70];
    assign x12_71 = in12[71];
    assign x12_72 = in12[72];
    wire x13_0;
    wire x13_1;
    wire x13_2;
    wire x13_3;
    wire x13_4;
    wire x13_5;
    wire x13_6;
    wire x13_7;
    wire x13_8;
    wire x13_9;
    wire x13_10;
    wire x13_11;
    wire x13_12;
    wire x13_13;
    wire x13_14;
    wire x13_15;
    wire x13_16;
    wire x13_17;
    wire x13_18;
    wire x13_19;
    wire x13_20;
    wire x13_21;
    wire x13_22;
    wire x13_23;
    wire x13_24;
    wire x13_25;
    wire x13_26;
    wire x13_27;
    wire x13_28;
    wire x13_29;
    wire x13_30;
    wire x13_31;
    wire x13_32;
    wire x13_33;
    wire x13_34;
    wire x13_35;
    wire x13_36;
    wire x13_37;
    wire x13_38;
    wire x13_39;
    wire x13_40;
    wire x13_41;
    wire x13_42;
    wire x13_43;
    wire x13_44;
    wire x13_45;
    wire x13_46;
    wire x13_47;
    wire x13_48;
    wire x13_49;
    wire x13_50;
    wire x13_51;
    wire x13_52;
    wire x13_53;
    wire x13_54;
    wire x13_55;
    wire x13_56;
    wire x13_57;
    wire x13_58;
    wire x13_59;
    wire x13_60;
    wire x13_61;
    wire x13_62;
    wire x13_63;
    wire x13_64;
    wire x13_65;
    wire x13_66;
    wire x13_67;
    wire x13_68;
    wire x13_69;
    wire x13_70;
    wire x13_71;
    wire x13_72;
    assign x13_0 = in13[0];
    assign x13_1 = in13[1];
    assign x13_2 = in13[2];
    assign x13_3 = in13[3];
    assign x13_4 = in13[4];
    assign x13_5 = in13[5];
    assign x13_6 = in13[6];
    assign x13_7 = in13[7];
    assign x13_8 = in13[8];
    assign x13_9 = in13[9];
    assign x13_10 = in13[10];
    assign x13_11 = in13[11];
    assign x13_12 = in13[12];
    assign x13_13 = in13[13];
    assign x13_14 = in13[14];
    assign x13_15 = in13[15];
    assign x13_16 = in13[16];
    assign x13_17 = in13[17];
    assign x13_18 = in13[18];
    assign x13_19 = in13[19];
    assign x13_20 = in13[20];
    assign x13_21 = in13[21];
    assign x13_22 = in13[22];
    assign x13_23 = in13[23];
    assign x13_24 = in13[24];
    assign x13_25 = in13[25];
    assign x13_26 = in13[26];
    assign x13_27 = in13[27];
    assign x13_28 = in13[28];
    assign x13_29 = in13[29];
    assign x13_30 = in13[30];
    assign x13_31 = in13[31];
    assign x13_32 = in13[32];
    assign x13_33 = in13[33];
    assign x13_34 = in13[34];
    assign x13_35 = in13[35];
    assign x13_36 = in13[36];
    assign x13_37 = in13[37];
    assign x13_38 = in13[38];
    assign x13_39 = in13[39];
    assign x13_40 = in13[40];
    assign x13_41 = in13[41];
    assign x13_42 = in13[42];
    assign x13_43 = in13[43];
    assign x13_44 = in13[44];
    assign x13_45 = in13[45];
    assign x13_46 = in13[46];
    assign x13_47 = in13[47];
    assign x13_48 = in13[48];
    assign x13_49 = in13[49];
    assign x13_50 = in13[50];
    assign x13_51 = in13[51];
    assign x13_52 = in13[52];
    assign x13_53 = in13[53];
    assign x13_54 = in13[54];
    assign x13_55 = in13[55];
    assign x13_56 = in13[56];
    assign x13_57 = in13[57];
    assign x13_58 = in13[58];
    assign x13_59 = in13[59];
    assign x13_60 = in13[60];
    assign x13_61 = in13[61];
    assign x13_62 = in13[62];
    assign x13_63 = in13[63];
    assign x13_64 = in13[64];
    assign x13_65 = in13[65];
    assign x13_66 = in13[66];
    assign x13_67 = in13[67];
    assign x13_68 = in13[68];
    assign x13_69 = in13[69];
    assign x13_70 = in13[70];
    assign x13_71 = in13[71];
    assign x13_72 = in13[72];
    wire x14_0;
    wire x14_1;
    wire x14_2;
    wire x14_3;
    wire x14_4;
    wire x14_5;
    wire x14_6;
    wire x14_7;
    wire x14_8;
    wire x14_9;
    wire x14_10;
    wire x14_11;
    wire x14_12;
    wire x14_13;
    wire x14_14;
    wire x14_15;
    wire x14_16;
    wire x14_17;
    wire x14_18;
    wire x14_19;
    wire x14_20;
    wire x14_21;
    wire x14_22;
    wire x14_23;
    wire x14_24;
    wire x14_25;
    wire x14_26;
    wire x14_27;
    wire x14_28;
    wire x14_29;
    wire x14_30;
    wire x14_31;
    wire x14_32;
    wire x14_33;
    wire x14_34;
    wire x14_35;
    wire x14_36;
    wire x14_37;
    wire x14_38;
    wire x14_39;
    wire x14_40;
    wire x14_41;
    wire x14_42;
    wire x14_43;
    wire x14_44;
    wire x14_45;
    wire x14_46;
    wire x14_47;
    wire x14_48;
    wire x14_49;
    wire x14_50;
    wire x14_51;
    wire x14_52;
    wire x14_53;
    wire x14_54;
    wire x14_55;
    wire x14_56;
    wire x14_57;
    wire x14_58;
    wire x14_59;
    wire x14_60;
    wire x14_61;
    wire x14_62;
    wire x14_63;
    wire x14_64;
    wire x14_65;
    wire x14_66;
    wire x14_67;
    wire x14_68;
    wire x14_69;
    wire x14_70;
    wire x14_71;
    wire x14_72;
    assign x14_0 = in14[0];
    assign x14_1 = in14[1];
    assign x14_2 = in14[2];
    assign x14_3 = in14[3];
    assign x14_4 = in14[4];
    assign x14_5 = in14[5];
    assign x14_6 = in14[6];
    assign x14_7 = in14[7];
    assign x14_8 = in14[8];
    assign x14_9 = in14[9];
    assign x14_10 = in14[10];
    assign x14_11 = in14[11];
    assign x14_12 = in14[12];
    assign x14_13 = in14[13];
    assign x14_14 = in14[14];
    assign x14_15 = in14[15];
    assign x14_16 = in14[16];
    assign x14_17 = in14[17];
    assign x14_18 = in14[18];
    assign x14_19 = in14[19];
    assign x14_20 = in14[20];
    assign x14_21 = in14[21];
    assign x14_22 = in14[22];
    assign x14_23 = in14[23];
    assign x14_24 = in14[24];
    assign x14_25 = in14[25];
    assign x14_26 = in14[26];
    assign x14_27 = in14[27];
    assign x14_28 = in14[28];
    assign x14_29 = in14[29];
    assign x14_30 = in14[30];
    assign x14_31 = in14[31];
    assign x14_32 = in14[32];
    assign x14_33 = in14[33];
    assign x14_34 = in14[34];
    assign x14_35 = in14[35];
    assign x14_36 = in14[36];
    assign x14_37 = in14[37];
    assign x14_38 = in14[38];
    assign x14_39 = in14[39];
    assign x14_40 = in14[40];
    assign x14_41 = in14[41];
    assign x14_42 = in14[42];
    assign x14_43 = in14[43];
    assign x14_44 = in14[44];
    assign x14_45 = in14[45];
    assign x14_46 = in14[46];
    assign x14_47 = in14[47];
    assign x14_48 = in14[48];
    assign x14_49 = in14[49];
    assign x14_50 = in14[50];
    assign x14_51 = in14[51];
    assign x14_52 = in14[52];
    assign x14_53 = in14[53];
    assign x14_54 = in14[54];
    assign x14_55 = in14[55];
    assign x14_56 = in14[56];
    assign x14_57 = in14[57];
    assign x14_58 = in14[58];
    assign x14_59 = in14[59];
    assign x14_60 = in14[60];
    assign x14_61 = in14[61];
    assign x14_62 = in14[62];
    assign x14_63 = in14[63];
    assign x14_64 = in14[64];
    assign x14_65 = in14[65];
    assign x14_66 = in14[66];
    assign x14_67 = in14[67];
    assign x14_68 = in14[68];
    assign x14_69 = in14[69];
    assign x14_70 = in14[70];
    assign x14_71 = in14[71];
    assign x14_72 = in14[72];
    wire x15_0;
    wire x15_1;
    wire x15_2;
    wire x15_3;
    wire x15_4;
    wire x15_5;
    wire x15_6;
    wire x15_7;
    wire x15_8;
    wire x15_9;
    wire x15_10;
    wire x15_11;
    wire x15_12;
    wire x15_13;
    wire x15_14;
    wire x15_15;
    wire x15_16;
    wire x15_17;
    wire x15_18;
    wire x15_19;
    wire x15_20;
    wire x15_21;
    wire x15_22;
    wire x15_23;
    wire x15_24;
    wire x15_25;
    wire x15_26;
    wire x15_27;
    wire x15_28;
    wire x15_29;
    wire x15_30;
    wire x15_31;
    wire x15_32;
    wire x15_33;
    wire x15_34;
    wire x15_35;
    wire x15_36;
    wire x15_37;
    wire x15_38;
    wire x15_39;
    wire x15_40;
    wire x15_41;
    wire x15_42;
    wire x15_43;
    wire x15_44;
    wire x15_45;
    wire x15_46;
    wire x15_47;
    wire x15_48;
    wire x15_49;
    wire x15_50;
    wire x15_51;
    wire x15_52;
    wire x15_53;
    wire x15_54;
    wire x15_55;
    wire x15_56;
    wire x15_57;
    wire x15_58;
    wire x15_59;
    wire x15_60;
    wire x15_61;
    wire x15_62;
    wire x15_63;
    wire x15_64;
    wire x15_65;
    wire x15_66;
    wire x15_67;
    wire x15_68;
    wire x15_69;
    wire x15_70;
    wire x15_71;
    wire x15_72;
    assign x15_0 = in15[0];
    assign x15_1 = in15[1];
    assign x15_2 = in15[2];
    assign x15_3 = in15[3];
    assign x15_4 = in15[4];
    assign x15_5 = in15[5];
    assign x15_6 = in15[6];
    assign x15_7 = in15[7];
    assign x15_8 = in15[8];
    assign x15_9 = in15[9];
    assign x15_10 = in15[10];
    assign x15_11 = in15[11];
    assign x15_12 = in15[12];
    assign x15_13 = in15[13];
    assign x15_14 = in15[14];
    assign x15_15 = in15[15];
    assign x15_16 = in15[16];
    assign x15_17 = in15[17];
    assign x15_18 = in15[18];
    assign x15_19 = in15[19];
    assign x15_20 = in15[20];
    assign x15_21 = in15[21];
    assign x15_22 = in15[22];
    assign x15_23 = in15[23];
    assign x15_24 = in15[24];
    assign x15_25 = in15[25];
    assign x15_26 = in15[26];
    assign x15_27 = in15[27];
    assign x15_28 = in15[28];
    assign x15_29 = in15[29];
    assign x15_30 = in15[30];
    assign x15_31 = in15[31];
    assign x15_32 = in15[32];
    assign x15_33 = in15[33];
    assign x15_34 = in15[34];
    assign x15_35 = in15[35];
    assign x15_36 = in15[36];
    assign x15_37 = in15[37];
    assign x15_38 = in15[38];
    assign x15_39 = in15[39];
    assign x15_40 = in15[40];
    assign x15_41 = in15[41];
    assign x15_42 = in15[42];
    assign x15_43 = in15[43];
    assign x15_44 = in15[44];
    assign x15_45 = in15[45];
    assign x15_46 = in15[46];
    assign x15_47 = in15[47];
    assign x15_48 = in15[48];
    assign x15_49 = in15[49];
    assign x15_50 = in15[50];
    assign x15_51 = in15[51];
    assign x15_52 = in15[52];
    assign x15_53 = in15[53];
    assign x15_54 = in15[54];
    assign x15_55 = in15[55];
    assign x15_56 = in15[56];
    assign x15_57 = in15[57];
    assign x15_58 = in15[58];
    assign x15_59 = in15[59];
    assign x15_60 = in15[60];
    assign x15_61 = in15[61];
    assign x15_62 = in15[62];
    assign x15_63 = in15[63];
    assign x15_64 = in15[64];
    assign x15_65 = in15[65];
    assign x15_66 = in15[66];
    assign x15_67 = in15[67];
    assign x15_68 = in15[68];
    assign x15_69 = in15[69];
    assign x15_70 = in15[70];
    assign x15_71 = in15[71];
    assign x15_72 = in15[72];
    wire w4688;
    wire w4689;
    wire w4690;
    wire w4691;
    wire w4692;
    wire w4693;
    wire w4694;
    wire w4695;
    wire w4696;
    wire w4697;
    wire w4698;
    wire w4699;
    wire w4700;
    wire w4701;
    wire w4702;
    wire w4703;
    wire w4704;
    wire w4705;
    wire w4706;
    wire w4707;
    wire w4708;
    wire w4709;
    wire w4710;
    wire w4711;
    wire w4712;
    wire w4713;
    wire w4714;
    wire w4715;
    wire w4716;
    wire w4717;
    wire w4718;
    wire w4719;
    wire w4720;
    wire w4721;
    wire w4722;
    wire w4723;
    wire w4724;
    wire w4725;
    wire w4726;
    wire w4727;
    wire w4728;
    wire w4729;
    wire w4730;
    wire w4731;
    wire w4732;
    wire w4733;
    wire w4734;
    wire w4735;
    wire w4736;
    wire w4737;
    wire w4738;
    wire w4739;
    wire w4740;
    wire w4741;
    wire w4742;
    wire w4743;
    wire w4744;
    wire w4745;
    wire w4746;
    wire w4747;
    wire w4748;
    wire w4749;
    wire w4750;
    wire w4751;
    wire w4752;
    wire w4753;
    wire w4754;
    wire w4755;
    wire w4756;
    wire w4761;
    wire w4762;
    wire w4763;
    wire w4764;
    assign out0[0] = w4688;
    assign out0[1] = w4689;
    assign out0[2] = w4690;
    assign out0[3] = w4691;
    assign out0[4] = w4692;
    assign out0[5] = w4693;
    assign out0[6] = w4694;
    assign out0[7] = w4695;
    assign out0[8] = w4696;
    assign out0[9] = w4697;
    assign out0[10] = w4698;
    assign out0[11] = w4699;
    assign out0[12] = w4700;
    assign out0[13] = w4701;
    assign out0[14] = w4702;
    assign out0[15] = w4703;
    assign out0[16] = w4704;
    assign out0[17] = w4705;
    assign out0[18] = w4706;
    assign out0[19] = w4707;
    assign out0[20] = w4708;
    assign out0[21] = w4709;
    assign out0[22] = w4710;
    assign out0[23] = w4711;
    assign out0[24] = w4712;
    assign out0[25] = w4713;
    assign out0[26] = w4714;
    assign out0[27] = w4715;
    assign out0[28] = w4716;
    assign out0[29] = w4717;
    assign out0[30] = w4718;
    assign out0[31] = w4719;
    assign out0[32] = w4720;
    assign out0[33] = w4721;
    assign out0[34] = w4722;
    assign out0[35] = w4723;
    assign out0[36] = w4724;
    assign out0[37] = w4725;
    assign out0[38] = w4726;
    assign out0[39] = w4727;
    assign out0[40] = w4728;
    assign out0[41] = w4729;
    assign out0[42] = w4730;
    assign out0[43] = w4731;
    assign out0[44] = w4732;
    assign out0[45] = w4733;
    assign out0[46] = w4734;
    assign out0[47] = w4735;
    assign out0[48] = w4736;
    assign out0[49] = w4737;
    assign out0[50] = w4738;
    assign out0[51] = w4739;
    assign out0[52] = w4740;
    assign out0[53] = w4741;
    assign out0[54] = w4742;
    assign out0[55] = w4743;
    assign out0[56] = w4744;
    assign out0[57] = w4745;
    assign out0[58] = w4746;
    assign out0[59] = w4747;
    assign out0[60] = w4748;
    assign out0[61] = w4749;
    assign out0[62] = w4750;
    assign out0[63] = w4751;
    assign out0[64] = w4752;
    assign out0[65] = w4753;
    assign out0[66] = w4754;
    assign out0[67] = w4755;
    assign out0[68] = w4756;
    assign out0[69] = w4761;
    assign out0[70] = w4762;
    assign out0[71] = w4763;
    assign out0[72] = w4764;
    wire w2909;
    wire w2910;
    wire w2911;
    wire w2912;
    wire w2913;
    wire w2914;
    wire w2915;
    wire w2916;
    wire w2917;
    wire w2918;
    wire w2919;
    wire w2920;
    wire w2921;
    wire w2922;
    wire w2923;
    wire w2924;
    wire w2925;
    wire w2926;
    wire w2927;
    wire w2928;
    wire w2929;
    wire w2930;
    wire w2931;
    wire w2932;
    wire w2933;
    wire w2934;
    wire w2935;
    wire w2936;
    wire w2937;
    wire w2938;
    wire w2939;
    wire w2940;
    wire w2941;
    wire w2942;
    wire w2943;
    wire w2944;
    wire w2945;
    wire w2946;
    wire w2947;
    wire w2948;
    wire w2949;
    wire w2950;
    wire w2951;
    wire w2952;
    wire w2953;
    wire w2954;
    wire w2955;
    wire w2956;
    wire w2957;
    wire w2958;
    wire w2959;
    wire w2960;
    wire w2961;
    wire w2962;
    wire w2963;
    wire w2964;
    wire w2965;
    wire w2966;
    wire w2967;
    wire w2968;
    wire w2969;
    wire w2970;
    wire w2971;
    wire w2972;
    wire w2973;
    wire w2974;
    wire w2975;
    wire w2976;
    wire w2977;
    wire w4765;
    wire w4766;
    wire w4767;
    wire w4768;
    assign out1[0] = w2909;
    assign out1[1] = w2910;
    assign out1[2] = w2911;
    assign out1[3] = w2912;
    assign out1[4] = w2913;
    assign out1[5] = w2914;
    assign out1[6] = w2915;
    assign out1[7] = w2916;
    assign out1[8] = w2917;
    assign out1[9] = w2918;
    assign out1[10] = w2919;
    assign out1[11] = w2920;
    assign out1[12] = w2921;
    assign out1[13] = w2922;
    assign out1[14] = w2923;
    assign out1[15] = w2924;
    assign out1[16] = w2925;
    assign out1[17] = w2926;
    assign out1[18] = w2927;
    assign out1[19] = w2928;
    assign out1[20] = w2929;
    assign out1[21] = w2930;
    assign out1[22] = w2931;
    assign out1[23] = w2932;
    assign out1[24] = w2933;
    assign out1[25] = w2934;
    assign out1[26] = w2935;
    assign out1[27] = w2936;
    assign out1[28] = w2937;
    assign out1[29] = w2938;
    assign out1[30] = w2939;
    assign out1[31] = w2940;
    assign out1[32] = w2941;
    assign out1[33] = w2942;
    assign out1[34] = w2943;
    assign out1[35] = w2944;
    assign out1[36] = w2945;
    assign out1[37] = w2946;
    assign out1[38] = w2947;
    assign out1[39] = w2948;
    assign out1[40] = w2949;
    assign out1[41] = w2950;
    assign out1[42] = w2951;
    assign out1[43] = w2952;
    assign out1[44] = w2953;
    assign out1[45] = w2954;
    assign out1[46] = w2955;
    assign out1[47] = w2956;
    assign out1[48] = w2957;
    assign out1[49] = w2958;
    assign out1[50] = w2959;
    assign out1[51] = w2960;
    assign out1[52] = w2961;
    assign out1[53] = w2962;
    assign out1[54] = w2963;
    assign out1[55] = w2964;
    assign out1[56] = w2965;
    assign out1[57] = w2966;
    assign out1[58] = w2967;
    assign out1[59] = w2968;
    assign out1[60] = w2969;
    assign out1[61] = w2970;
    assign out1[62] = w2971;
    assign out1[63] = w2972;
    assign out1[64] = w2973;
    assign out1[65] = w2974;
    assign out1[66] = w2975;
    assign out1[67] = w2976;
    assign out1[68] = w2977;
    assign out1[69] = w4765;
    assign out1[70] = w4766;
    assign out1[71] = w4767;
    assign out1[72] = w4768;
    wire w4098;
    wire w4099;
    wire w4100;
    wire w4101;
    wire w4102;
    wire w4103;
    wire w4104;
    wire w4105;
    wire w4106;
    wire w4107;
    wire w4108;
    wire w4109;
    wire w4110;
    wire w4111;
    wire w4112;
    wire w4113;
    wire w4114;
    wire w4115;
    wire w4116;
    wire w4117;
    wire w4118;
    wire w4119;
    wire w4120;
    wire w4121;
    wire w4122;
    wire w4123;
    wire w4124;
    wire w4125;
    wire w4126;
    wire w4127;
    wire w4128;
    wire w4129;
    wire w4130;
    wire w4131;
    wire w4132;
    wire w4133;
    wire w4134;
    wire w4135;
    wire w4136;
    wire w4137;
    wire w4138;
    wire w4139;
    wire w4140;
    wire w4141;
    wire w4142;
    wire w4143;
    wire w4144;
    wire w4145;
    wire w4146;
    wire w4147;
    wire w4148;
    wire w4149;
    wire w4150;
    wire w4151;
    wire w4152;
    wire w4153;
    wire w4154;
    wire w4155;
    wire w4156;
    wire w4157;
    wire w4158;
    wire w4159;
    wire w4160;
    wire w4161;
    wire w4162;
    wire w4163;
    wire w4164;
    wire w4165;
    wire w4166;
    wire w4769;
    wire w4770;
    wire w4771;
    wire w4772;
    assign out2[0] = w4098;
    assign out2[1] = w4099;
    assign out2[2] = w4100;
    assign out2[3] = w4101;
    assign out2[4] = w4102;
    assign out2[5] = w4103;
    assign out2[6] = w4104;
    assign out2[7] = w4105;
    assign out2[8] = w4106;
    assign out2[9] = w4107;
    assign out2[10] = w4108;
    assign out2[11] = w4109;
    assign out2[12] = w4110;
    assign out2[13] = w4111;
    assign out2[14] = w4112;
    assign out2[15] = w4113;
    assign out2[16] = w4114;
    assign out2[17] = w4115;
    assign out2[18] = w4116;
    assign out2[19] = w4117;
    assign out2[20] = w4118;
    assign out2[21] = w4119;
    assign out2[22] = w4120;
    assign out2[23] = w4121;
    assign out2[24] = w4122;
    assign out2[25] = w4123;
    assign out2[26] = w4124;
    assign out2[27] = w4125;
    assign out2[28] = w4126;
    assign out2[29] = w4127;
    assign out2[30] = w4128;
    assign out2[31] = w4129;
    assign out2[32] = w4130;
    assign out2[33] = w4131;
    assign out2[34] = w4132;
    assign out2[35] = w4133;
    assign out2[36] = w4134;
    assign out2[37] = w4135;
    assign out2[38] = w4136;
    assign out2[39] = w4137;
    assign out2[40] = w4138;
    assign out2[41] = w4139;
    assign out2[42] = w4140;
    assign out2[43] = w4141;
    assign out2[44] = w4142;
    assign out2[45] = w4143;
    assign out2[46] = w4144;
    assign out2[47] = w4145;
    assign out2[48] = w4146;
    assign out2[49] = w4147;
    assign out2[50] = w4148;
    assign out2[51] = w4149;
    assign out2[52] = w4150;
    assign out2[53] = w4151;
    assign out2[54] = w4152;
    assign out2[55] = w4153;
    assign out2[56] = w4154;
    assign out2[57] = w4155;
    assign out2[58] = w4156;
    assign out2[59] = w4157;
    assign out2[60] = w4158;
    assign out2[61] = w4159;
    assign out2[62] = w4160;
    assign out2[63] = w4161;
    assign out2[64] = w4162;
    assign out2[65] = w4163;
    assign out2[66] = w4164;
    assign out2[67] = w4165;
    assign out2[68] = w4166;
    assign out2[69] = w4769;
    assign out2[70] = w4770;
    assign out2[71] = w4771;
    assign out2[72] = w4772;
    wire w2319;
    wire w2320;
    wire w2321;
    wire w2322;
    wire w2323;
    wire w2324;
    wire w2325;
    wire w2326;
    wire w2327;
    wire w2328;
    wire w2329;
    wire w2330;
    wire w2331;
    wire w2332;
    wire w2333;
    wire w2334;
    wire w2335;
    wire w2336;
    wire w2337;
    wire w2338;
    wire w2339;
    wire w2340;
    wire w2341;
    wire w2342;
    wire w2343;
    wire w2344;
    wire w2345;
    wire w2346;
    wire w2347;
    wire w2348;
    wire w2349;
    wire w2350;
    wire w2351;
    wire w2352;
    wire w2353;
    wire w2354;
    wire w2355;
    wire w2356;
    wire w2357;
    wire w2358;
    wire w2359;
    wire w2360;
    wire w2361;
    wire w2362;
    wire w2363;
    wire w2364;
    wire w2365;
    wire w2366;
    wire w2367;
    wire w2368;
    wire w2369;
    wire w2370;
    wire w2371;
    wire w2372;
    wire w2373;
    wire w2374;
    wire w2375;
    wire w2376;
    wire w2377;
    wire w2378;
    wire w2379;
    wire w2380;
    wire w2381;
    wire w2382;
    wire w2383;
    wire w2384;
    wire w2385;
    wire w2386;
    wire w2387;
    wire w4773;
    wire w4774;
    wire w4775;
    wire w4776;
    assign out3[0] = w2319;
    assign out3[1] = w2320;
    assign out3[2] = w2321;
    assign out3[3] = w2322;
    assign out3[4] = w2323;
    assign out3[5] = w2324;
    assign out3[6] = w2325;
    assign out3[7] = w2326;
    assign out3[8] = w2327;
    assign out3[9] = w2328;
    assign out3[10] = w2329;
    assign out3[11] = w2330;
    assign out3[12] = w2331;
    assign out3[13] = w2332;
    assign out3[14] = w2333;
    assign out3[15] = w2334;
    assign out3[16] = w2335;
    assign out3[17] = w2336;
    assign out3[18] = w2337;
    assign out3[19] = w2338;
    assign out3[20] = w2339;
    assign out3[21] = w2340;
    assign out3[22] = w2341;
    assign out3[23] = w2342;
    assign out3[24] = w2343;
    assign out3[25] = w2344;
    assign out3[26] = w2345;
    assign out3[27] = w2346;
    assign out3[28] = w2347;
    assign out3[29] = w2348;
    assign out3[30] = w2349;
    assign out3[31] = w2350;
    assign out3[32] = w2351;
    assign out3[33] = w2352;
    assign out3[34] = w2353;
    assign out3[35] = w2354;
    assign out3[36] = w2355;
    assign out3[37] = w2356;
    assign out3[38] = w2357;
    assign out3[39] = w2358;
    assign out3[40] = w2359;
    assign out3[41] = w2360;
    assign out3[42] = w2361;
    assign out3[43] = w2362;
    assign out3[44] = w2363;
    assign out3[45] = w2364;
    assign out3[46] = w2365;
    assign out3[47] = w2366;
    assign out3[48] = w2367;
    assign out3[49] = w2368;
    assign out3[50] = w2369;
    assign out3[51] = w2370;
    assign out3[52] = w2371;
    assign out3[53] = w2372;
    assign out3[54] = w2373;
    assign out3[55] = w2374;
    assign out3[56] = w2375;
    assign out3[57] = w2376;
    assign out3[58] = w2377;
    assign out3[59] = w2378;
    assign out3[60] = w2379;
    assign out3[61] = w2380;
    assign out3[62] = w2381;
    assign out3[63] = w2382;
    assign out3[64] = w2383;
    assign out3[65] = w2384;
    assign out3[66] = w2385;
    assign out3[67] = w2386;
    assign out3[68] = w2387;
    assign out3[69] = w4773;
    assign out3[70] = w4774;
    assign out3[71] = w4775;
    assign out3[72] = w4776;
    wire w4542;
    wire w4543;
    wire w4544;
    wire w4545;
    wire w4546;
    wire w4547;
    wire w4548;
    wire w4549;
    wire w4550;
    wire w4551;
    wire w4552;
    wire w4553;
    wire w4554;
    wire w4555;
    wire w4556;
    wire w4557;
    wire w4558;
    wire w4559;
    wire w4560;
    wire w4561;
    wire w4562;
    wire w4563;
    wire w4564;
    wire w4565;
    wire w4566;
    wire w4567;
    wire w4568;
    wire w4569;
    wire w4570;
    wire w4571;
    wire w4572;
    wire w4573;
    wire w4574;
    wire w4575;
    wire w4576;
    wire w4577;
    wire w4578;
    wire w4579;
    wire w4580;
    wire w4581;
    wire w4582;
    wire w4583;
    wire w4584;
    wire w4585;
    wire w4586;
    wire w4587;
    wire w4588;
    wire w4589;
    wire w4590;
    wire w4591;
    wire w4592;
    wire w4593;
    wire w4594;
    wire w4595;
    wire w4596;
    wire w4597;
    wire w4598;
    wire w4599;
    wire w4600;
    wire w4601;
    wire w4602;
    wire w4603;
    wire w4604;
    wire w4605;
    wire w4606;
    wire w4607;
    wire w4608;
    wire w4609;
    wire w4610;
    wire w4777;
    wire w4778;
    wire w4779;
    wire w4780;
    assign out4[0] = w4542;
    assign out4[1] = w4543;
    assign out4[2] = w4544;
    assign out4[3] = w4545;
    assign out4[4] = w4546;
    assign out4[5] = w4547;
    assign out4[6] = w4548;
    assign out4[7] = w4549;
    assign out4[8] = w4550;
    assign out4[9] = w4551;
    assign out4[10] = w4552;
    assign out4[11] = w4553;
    assign out4[12] = w4554;
    assign out4[13] = w4555;
    assign out4[14] = w4556;
    assign out4[15] = w4557;
    assign out4[16] = w4558;
    assign out4[17] = w4559;
    assign out4[18] = w4560;
    assign out4[19] = w4561;
    assign out4[20] = w4562;
    assign out4[21] = w4563;
    assign out4[22] = w4564;
    assign out4[23] = w4565;
    assign out4[24] = w4566;
    assign out4[25] = w4567;
    assign out4[26] = w4568;
    assign out4[27] = w4569;
    assign out4[28] = w4570;
    assign out4[29] = w4571;
    assign out4[30] = w4572;
    assign out4[31] = w4573;
    assign out4[32] = w4574;
    assign out4[33] = w4575;
    assign out4[34] = w4576;
    assign out4[35] = w4577;
    assign out4[36] = w4578;
    assign out4[37] = w4579;
    assign out4[38] = w4580;
    assign out4[39] = w4581;
    assign out4[40] = w4582;
    assign out4[41] = w4583;
    assign out4[42] = w4584;
    assign out4[43] = w4585;
    assign out4[44] = w4586;
    assign out4[45] = w4587;
    assign out4[46] = w4588;
    assign out4[47] = w4589;
    assign out4[48] = w4590;
    assign out4[49] = w4591;
    assign out4[50] = w4592;
    assign out4[51] = w4593;
    assign out4[52] = w4594;
    assign out4[53] = w4595;
    assign out4[54] = w4596;
    assign out4[55] = w4597;
    assign out4[56] = w4598;
    assign out4[57] = w4599;
    assign out4[58] = w4600;
    assign out4[59] = w4601;
    assign out4[60] = w4602;
    assign out4[61] = w4603;
    assign out4[62] = w4604;
    assign out4[63] = w4605;
    assign out4[64] = w4606;
    assign out4[65] = w4607;
    assign out4[66] = w4608;
    assign out4[67] = w4609;
    assign out4[68] = w4610;
    assign out4[69] = w4777;
    assign out4[70] = w4778;
    assign out4[71] = w4779;
    assign out4[72] = w4780;
    wire w2763;
    wire w2764;
    wire w2765;
    wire w2766;
    wire w2767;
    wire w2768;
    wire w2769;
    wire w2770;
    wire w2771;
    wire w2772;
    wire w2773;
    wire w2774;
    wire w2775;
    wire w2776;
    wire w2777;
    wire w2778;
    wire w2779;
    wire w2780;
    wire w2781;
    wire w2782;
    wire w2783;
    wire w2784;
    wire w2785;
    wire w2786;
    wire w2787;
    wire w2788;
    wire w2789;
    wire w2790;
    wire w2791;
    wire w2792;
    wire w2793;
    wire w2794;
    wire w2795;
    wire w2796;
    wire w2797;
    wire w2798;
    wire w2799;
    wire w2800;
    wire w2801;
    wire w2802;
    wire w2803;
    wire w2804;
    wire w2805;
    wire w2806;
    wire w2807;
    wire w2808;
    wire w2809;
    wire w2810;
    wire w2811;
    wire w2812;
    wire w2813;
    wire w2814;
    wire w2815;
    wire w2816;
    wire w2817;
    wire w2818;
    wire w2819;
    wire w2820;
    wire w2821;
    wire w2822;
    wire w2823;
    wire w2824;
    wire w2825;
    wire w2826;
    wire w2827;
    wire w2828;
    wire w2829;
    wire w2830;
    wire w2831;
    wire w4781;
    wire w4782;
    wire w4783;
    wire w4784;
    assign out5[0] = w2763;
    assign out5[1] = w2764;
    assign out5[2] = w2765;
    assign out5[3] = w2766;
    assign out5[4] = w2767;
    assign out5[5] = w2768;
    assign out5[6] = w2769;
    assign out5[7] = w2770;
    assign out5[8] = w2771;
    assign out5[9] = w2772;
    assign out5[10] = w2773;
    assign out5[11] = w2774;
    assign out5[12] = w2775;
    assign out5[13] = w2776;
    assign out5[14] = w2777;
    assign out5[15] = w2778;
    assign out5[16] = w2779;
    assign out5[17] = w2780;
    assign out5[18] = w2781;
    assign out5[19] = w2782;
    assign out5[20] = w2783;
    assign out5[21] = w2784;
    assign out5[22] = w2785;
    assign out5[23] = w2786;
    assign out5[24] = w2787;
    assign out5[25] = w2788;
    assign out5[26] = w2789;
    assign out5[27] = w2790;
    assign out5[28] = w2791;
    assign out5[29] = w2792;
    assign out5[30] = w2793;
    assign out5[31] = w2794;
    assign out5[32] = w2795;
    assign out5[33] = w2796;
    assign out5[34] = w2797;
    assign out5[35] = w2798;
    assign out5[36] = w2799;
    assign out5[37] = w2800;
    assign out5[38] = w2801;
    assign out5[39] = w2802;
    assign out5[40] = w2803;
    assign out5[41] = w2804;
    assign out5[42] = w2805;
    assign out5[43] = w2806;
    assign out5[44] = w2807;
    assign out5[45] = w2808;
    assign out5[46] = w2809;
    assign out5[47] = w2810;
    assign out5[48] = w2811;
    assign out5[49] = w2812;
    assign out5[50] = w2813;
    assign out5[51] = w2814;
    assign out5[52] = w2815;
    assign out5[53] = w2816;
    assign out5[54] = w2817;
    assign out5[55] = w2818;
    assign out5[56] = w2819;
    assign out5[57] = w2820;
    assign out5[58] = w2821;
    assign out5[59] = w2822;
    assign out5[60] = w2823;
    assign out5[61] = w2824;
    assign out5[62] = w2825;
    assign out5[63] = w2826;
    assign out5[64] = w2827;
    assign out5[65] = w2828;
    assign out5[66] = w2829;
    assign out5[67] = w2830;
    assign out5[68] = w2831;
    assign out5[69] = w4781;
    assign out5[70] = w4782;
    assign out5[71] = w4783;
    assign out5[72] = w4784;
    wire w3952;
    wire w3953;
    wire w3954;
    wire w3955;
    wire w3956;
    wire w3957;
    wire w3958;
    wire w3959;
    wire w3960;
    wire w3961;
    wire w3962;
    wire w3963;
    wire w3964;
    wire w3965;
    wire w3966;
    wire w3967;
    wire w3968;
    wire w3969;
    wire w3970;
    wire w3971;
    wire w3972;
    wire w3973;
    wire w3974;
    wire w3975;
    wire w3976;
    wire w3977;
    wire w3978;
    wire w3979;
    wire w3980;
    wire w3981;
    wire w3982;
    wire w3983;
    wire w3984;
    wire w3985;
    wire w3986;
    wire w3987;
    wire w3988;
    wire w3989;
    wire w3990;
    wire w3991;
    wire w3992;
    wire w3993;
    wire w3994;
    wire w3995;
    wire w3996;
    wire w3997;
    wire w3998;
    wire w3999;
    wire w4000;
    wire w4001;
    wire w4002;
    wire w4003;
    wire w4004;
    wire w4005;
    wire w4006;
    wire w4007;
    wire w4008;
    wire w4009;
    wire w4010;
    wire w4011;
    wire w4012;
    wire w4013;
    wire w4014;
    wire w4015;
    wire w4016;
    wire w4017;
    wire w4018;
    wire w4019;
    wire w4020;
    wire w4785;
    wire w4786;
    wire w4787;
    wire w4788;
    assign out6[0] = w3952;
    assign out6[1] = w3953;
    assign out6[2] = w3954;
    assign out6[3] = w3955;
    assign out6[4] = w3956;
    assign out6[5] = w3957;
    assign out6[6] = w3958;
    assign out6[7] = w3959;
    assign out6[8] = w3960;
    assign out6[9] = w3961;
    assign out6[10] = w3962;
    assign out6[11] = w3963;
    assign out6[12] = w3964;
    assign out6[13] = w3965;
    assign out6[14] = w3966;
    assign out6[15] = w3967;
    assign out6[16] = w3968;
    assign out6[17] = w3969;
    assign out6[18] = w3970;
    assign out6[19] = w3971;
    assign out6[20] = w3972;
    assign out6[21] = w3973;
    assign out6[22] = w3974;
    assign out6[23] = w3975;
    assign out6[24] = w3976;
    assign out6[25] = w3977;
    assign out6[26] = w3978;
    assign out6[27] = w3979;
    assign out6[28] = w3980;
    assign out6[29] = w3981;
    assign out6[30] = w3982;
    assign out6[31] = w3983;
    assign out6[32] = w3984;
    assign out6[33] = w3985;
    assign out6[34] = w3986;
    assign out6[35] = w3987;
    assign out6[36] = w3988;
    assign out6[37] = w3989;
    assign out6[38] = w3990;
    assign out6[39] = w3991;
    assign out6[40] = w3992;
    assign out6[41] = w3993;
    assign out6[42] = w3994;
    assign out6[43] = w3995;
    assign out6[44] = w3996;
    assign out6[45] = w3997;
    assign out6[46] = w3998;
    assign out6[47] = w3999;
    assign out6[48] = w4000;
    assign out6[49] = w4001;
    assign out6[50] = w4002;
    assign out6[51] = w4003;
    assign out6[52] = w4004;
    assign out6[53] = w4005;
    assign out6[54] = w4006;
    assign out6[55] = w4007;
    assign out6[56] = w4008;
    assign out6[57] = w4009;
    assign out6[58] = w4010;
    assign out6[59] = w4011;
    assign out6[60] = w4012;
    assign out6[61] = w4013;
    assign out6[62] = w4014;
    assign out6[63] = w4015;
    assign out6[64] = w4016;
    assign out6[65] = w4017;
    assign out6[66] = w4018;
    assign out6[67] = w4019;
    assign out6[68] = w4020;
    assign out6[69] = w4785;
    assign out6[70] = w4786;
    assign out6[71] = w4787;
    assign out6[72] = w4788;
    wire w2173;
    wire w2174;
    wire w2175;
    wire w2176;
    wire w2177;
    wire w2178;
    wire w2179;
    wire w2180;
    wire w2181;
    wire w2182;
    wire w2183;
    wire w2184;
    wire w2185;
    wire w2186;
    wire w2187;
    wire w2188;
    wire w2189;
    wire w2190;
    wire w2191;
    wire w2192;
    wire w2193;
    wire w2194;
    wire w2195;
    wire w2196;
    wire w2197;
    wire w2198;
    wire w2199;
    wire w2200;
    wire w2201;
    wire w2202;
    wire w2203;
    wire w2204;
    wire w2205;
    wire w2206;
    wire w2207;
    wire w2208;
    wire w2209;
    wire w2210;
    wire w2211;
    wire w2212;
    wire w2213;
    wire w2214;
    wire w2215;
    wire w2216;
    wire w2217;
    wire w2218;
    wire w2219;
    wire w2220;
    wire w2221;
    wire w2222;
    wire w2223;
    wire w2224;
    wire w2225;
    wire w2226;
    wire w2227;
    wire w2228;
    wire w2229;
    wire w2230;
    wire w2231;
    wire w2232;
    wire w2233;
    wire w2234;
    wire w2235;
    wire w2236;
    wire w2237;
    wire w2238;
    wire w2239;
    wire w2240;
    wire w2241;
    wire w4789;
    wire w4790;
    wire w4791;
    wire w4792;
    assign out7[0] = w2173;
    assign out7[1] = w2174;
    assign out7[2] = w2175;
    assign out7[3] = w2176;
    assign out7[4] = w2177;
    assign out7[5] = w2178;
    assign out7[6] = w2179;
    assign out7[7] = w2180;
    assign out7[8] = w2181;
    assign out7[9] = w2182;
    assign out7[10] = w2183;
    assign out7[11] = w2184;
    assign out7[12] = w2185;
    assign out7[13] = w2186;
    assign out7[14] = w2187;
    assign out7[15] = w2188;
    assign out7[16] = w2189;
    assign out7[17] = w2190;
    assign out7[18] = w2191;
    assign out7[19] = w2192;
    assign out7[20] = w2193;
    assign out7[21] = w2194;
    assign out7[22] = w2195;
    assign out7[23] = w2196;
    assign out7[24] = w2197;
    assign out7[25] = w2198;
    assign out7[26] = w2199;
    assign out7[27] = w2200;
    assign out7[28] = w2201;
    assign out7[29] = w2202;
    assign out7[30] = w2203;
    assign out7[31] = w2204;
    assign out7[32] = w2205;
    assign out7[33] = w2206;
    assign out7[34] = w2207;
    assign out7[35] = w2208;
    assign out7[36] = w2209;
    assign out7[37] = w2210;
    assign out7[38] = w2211;
    assign out7[39] = w2212;
    assign out7[40] = w2213;
    assign out7[41] = w2214;
    assign out7[42] = w2215;
    assign out7[43] = w2216;
    assign out7[44] = w2217;
    assign out7[45] = w2218;
    assign out7[46] = w2219;
    assign out7[47] = w2220;
    assign out7[48] = w2221;
    assign out7[49] = w2222;
    assign out7[50] = w2223;
    assign out7[51] = w2224;
    assign out7[52] = w2225;
    assign out7[53] = w2226;
    assign out7[54] = w2227;
    assign out7[55] = w2228;
    assign out7[56] = w2229;
    assign out7[57] = w2230;
    assign out7[58] = w2231;
    assign out7[59] = w2232;
    assign out7[60] = w2233;
    assign out7[61] = w2234;
    assign out7[62] = w2235;
    assign out7[63] = w2236;
    assign out7[64] = w2237;
    assign out7[65] = w2238;
    assign out7[66] = w2239;
    assign out7[67] = w2240;
    assign out7[68] = w2241;
    assign out7[69] = w4789;
    assign out7[70] = w4790;
    assign out7[71] = w4791;
    assign out7[72] = w4792;
    wire w4615;
    wire w4616;
    wire w4617;
    wire w4618;
    wire w4619;
    wire w4620;
    wire w4621;
    wire w4622;
    wire w4623;
    wire w4624;
    wire w4625;
    wire w4626;
    wire w4627;
    wire w4628;
    wire w4629;
    wire w4630;
    wire w4631;
    wire w4632;
    wire w4633;
    wire w4634;
    wire w4635;
    wire w4636;
    wire w4637;
    wire w4638;
    wire w4639;
    wire w4640;
    wire w4641;
    wire w4642;
    wire w4643;
    wire w4644;
    wire w4645;
    wire w4646;
    wire w4647;
    wire w4648;
    wire w4649;
    wire w4650;
    wire w4651;
    wire w4652;
    wire w4653;
    wire w4654;
    wire w4655;
    wire w4656;
    wire w4657;
    wire w4658;
    wire w4659;
    wire w4660;
    wire w4661;
    wire w4662;
    wire w4663;
    wire w4664;
    wire w4665;
    wire w4666;
    wire w4667;
    wire w4668;
    wire w4669;
    wire w4670;
    wire w4671;
    wire w4672;
    wire w4673;
    wire w4674;
    wire w4675;
    wire w4676;
    wire w4677;
    wire w4678;
    wire w4679;
    wire w4680;
    wire w4681;
    wire w4682;
    wire w4683;
    wire w4793;
    wire w4794;
    wire w4795;
    wire w4796;
    assign out8[0] = w4615;
    assign out8[1] = w4616;
    assign out8[2] = w4617;
    assign out8[3] = w4618;
    assign out8[4] = w4619;
    assign out8[5] = w4620;
    assign out8[6] = w4621;
    assign out8[7] = w4622;
    assign out8[8] = w4623;
    assign out8[9] = w4624;
    assign out8[10] = w4625;
    assign out8[11] = w4626;
    assign out8[12] = w4627;
    assign out8[13] = w4628;
    assign out8[14] = w4629;
    assign out8[15] = w4630;
    assign out8[16] = w4631;
    assign out8[17] = w4632;
    assign out8[18] = w4633;
    assign out8[19] = w4634;
    assign out8[20] = w4635;
    assign out8[21] = w4636;
    assign out8[22] = w4637;
    assign out8[23] = w4638;
    assign out8[24] = w4639;
    assign out8[25] = w4640;
    assign out8[26] = w4641;
    assign out8[27] = w4642;
    assign out8[28] = w4643;
    assign out8[29] = w4644;
    assign out8[30] = w4645;
    assign out8[31] = w4646;
    assign out8[32] = w4647;
    assign out8[33] = w4648;
    assign out8[34] = w4649;
    assign out8[35] = w4650;
    assign out8[36] = w4651;
    assign out8[37] = w4652;
    assign out8[38] = w4653;
    assign out8[39] = w4654;
    assign out8[40] = w4655;
    assign out8[41] = w4656;
    assign out8[42] = w4657;
    assign out8[43] = w4658;
    assign out8[44] = w4659;
    assign out8[45] = w4660;
    assign out8[46] = w4661;
    assign out8[47] = w4662;
    assign out8[48] = w4663;
    assign out8[49] = w4664;
    assign out8[50] = w4665;
    assign out8[51] = w4666;
    assign out8[52] = w4667;
    assign out8[53] = w4668;
    assign out8[54] = w4669;
    assign out8[55] = w4670;
    assign out8[56] = w4671;
    assign out8[57] = w4672;
    assign out8[58] = w4673;
    assign out8[59] = w4674;
    assign out8[60] = w4675;
    assign out8[61] = w4676;
    assign out8[62] = w4677;
    assign out8[63] = w4678;
    assign out8[64] = w4679;
    assign out8[65] = w4680;
    assign out8[66] = w4681;
    assign out8[67] = w4682;
    assign out8[68] = w4683;
    assign out8[69] = w4793;
    assign out8[70] = w4794;
    assign out8[71] = w4795;
    assign out8[72] = w4796;
    wire w2836;
    wire w2837;
    wire w2838;
    wire w2839;
    wire w2840;
    wire w2841;
    wire w2842;
    wire w2843;
    wire w2844;
    wire w2845;
    wire w2846;
    wire w2847;
    wire w2848;
    wire w2849;
    wire w2850;
    wire w2851;
    wire w2852;
    wire w2853;
    wire w2854;
    wire w2855;
    wire w2856;
    wire w2857;
    wire w2858;
    wire w2859;
    wire w2860;
    wire w2861;
    wire w2862;
    wire w2863;
    wire w2864;
    wire w2865;
    wire w2866;
    wire w2867;
    wire w2868;
    wire w2869;
    wire w2870;
    wire w2871;
    wire w2872;
    wire w2873;
    wire w2874;
    wire w2875;
    wire w2876;
    wire w2877;
    wire w2878;
    wire w2879;
    wire w2880;
    wire w2881;
    wire w2882;
    wire w2883;
    wire w2884;
    wire w2885;
    wire w2886;
    wire w2887;
    wire w2888;
    wire w2889;
    wire w2890;
    wire w2891;
    wire w2892;
    wire w2893;
    wire w2894;
    wire w2895;
    wire w2896;
    wire w2897;
    wire w2898;
    wire w2899;
    wire w2900;
    wire w2901;
    wire w2902;
    wire w2903;
    wire w2904;
    wire w4797;
    wire w4798;
    wire w4799;
    wire w4800;
    assign out9[0] = w2836;
    assign out9[1] = w2837;
    assign out9[2] = w2838;
    assign out9[3] = w2839;
    assign out9[4] = w2840;
    assign out9[5] = w2841;
    assign out9[6] = w2842;
    assign out9[7] = w2843;
    assign out9[8] = w2844;
    assign out9[9] = w2845;
    assign out9[10] = w2846;
    assign out9[11] = w2847;
    assign out9[12] = w2848;
    assign out9[13] = w2849;
    assign out9[14] = w2850;
    assign out9[15] = w2851;
    assign out9[16] = w2852;
    assign out9[17] = w2853;
    assign out9[18] = w2854;
    assign out9[19] = w2855;
    assign out9[20] = w2856;
    assign out9[21] = w2857;
    assign out9[22] = w2858;
    assign out9[23] = w2859;
    assign out9[24] = w2860;
    assign out9[25] = w2861;
    assign out9[26] = w2862;
    assign out9[27] = w2863;
    assign out9[28] = w2864;
    assign out9[29] = w2865;
    assign out9[30] = w2866;
    assign out9[31] = w2867;
    assign out9[32] = w2868;
    assign out9[33] = w2869;
    assign out9[34] = w2870;
    assign out9[35] = w2871;
    assign out9[36] = w2872;
    assign out9[37] = w2873;
    assign out9[38] = w2874;
    assign out9[39] = w2875;
    assign out9[40] = w2876;
    assign out9[41] = w2877;
    assign out9[42] = w2878;
    assign out9[43] = w2879;
    assign out9[44] = w2880;
    assign out9[45] = w2881;
    assign out9[46] = w2882;
    assign out9[47] = w2883;
    assign out9[48] = w2884;
    assign out9[49] = w2885;
    assign out9[50] = w2886;
    assign out9[51] = w2887;
    assign out9[52] = w2888;
    assign out9[53] = w2889;
    assign out9[54] = w2890;
    assign out9[55] = w2891;
    assign out9[56] = w2892;
    assign out9[57] = w2893;
    assign out9[58] = w2894;
    assign out9[59] = w2895;
    assign out9[60] = w2896;
    assign out9[61] = w2897;
    assign out9[62] = w2898;
    assign out9[63] = w2899;
    assign out9[64] = w2900;
    assign out9[65] = w2901;
    assign out9[66] = w2902;
    assign out9[67] = w2903;
    assign out9[68] = w2904;
    assign out9[69] = w4797;
    assign out9[70] = w4798;
    assign out9[71] = w4799;
    assign out9[72] = w4800;
    wire w4025;
    wire w4026;
    wire w4027;
    wire w4028;
    wire w4029;
    wire w4030;
    wire w4031;
    wire w4032;
    wire w4033;
    wire w4034;
    wire w4035;
    wire w4036;
    wire w4037;
    wire w4038;
    wire w4039;
    wire w4040;
    wire w4041;
    wire w4042;
    wire w4043;
    wire w4044;
    wire w4045;
    wire w4046;
    wire w4047;
    wire w4048;
    wire w4049;
    wire w4050;
    wire w4051;
    wire w4052;
    wire w4053;
    wire w4054;
    wire w4055;
    wire w4056;
    wire w4057;
    wire w4058;
    wire w4059;
    wire w4060;
    wire w4061;
    wire w4062;
    wire w4063;
    wire w4064;
    wire w4065;
    wire w4066;
    wire w4067;
    wire w4068;
    wire w4069;
    wire w4070;
    wire w4071;
    wire w4072;
    wire w4073;
    wire w4074;
    wire w4075;
    wire w4076;
    wire w4077;
    wire w4078;
    wire w4079;
    wire w4080;
    wire w4081;
    wire w4082;
    wire w4083;
    wire w4084;
    wire w4085;
    wire w4086;
    wire w4087;
    wire w4088;
    wire w4089;
    wire w4090;
    wire w4091;
    wire w4092;
    wire w4093;
    wire w4801;
    wire w4802;
    wire w4803;
    wire w4804;
    assign out10[0] = w4025;
    assign out10[1] = w4026;
    assign out10[2] = w4027;
    assign out10[3] = w4028;
    assign out10[4] = w4029;
    assign out10[5] = w4030;
    assign out10[6] = w4031;
    assign out10[7] = w4032;
    assign out10[8] = w4033;
    assign out10[9] = w4034;
    assign out10[10] = w4035;
    assign out10[11] = w4036;
    assign out10[12] = w4037;
    assign out10[13] = w4038;
    assign out10[14] = w4039;
    assign out10[15] = w4040;
    assign out10[16] = w4041;
    assign out10[17] = w4042;
    assign out10[18] = w4043;
    assign out10[19] = w4044;
    assign out10[20] = w4045;
    assign out10[21] = w4046;
    assign out10[22] = w4047;
    assign out10[23] = w4048;
    assign out10[24] = w4049;
    assign out10[25] = w4050;
    assign out10[26] = w4051;
    assign out10[27] = w4052;
    assign out10[28] = w4053;
    assign out10[29] = w4054;
    assign out10[30] = w4055;
    assign out10[31] = w4056;
    assign out10[32] = w4057;
    assign out10[33] = w4058;
    assign out10[34] = w4059;
    assign out10[35] = w4060;
    assign out10[36] = w4061;
    assign out10[37] = w4062;
    assign out10[38] = w4063;
    assign out10[39] = w4064;
    assign out10[40] = w4065;
    assign out10[41] = w4066;
    assign out10[42] = w4067;
    assign out10[43] = w4068;
    assign out10[44] = w4069;
    assign out10[45] = w4070;
    assign out10[46] = w4071;
    assign out10[47] = w4072;
    assign out10[48] = w4073;
    assign out10[49] = w4074;
    assign out10[50] = w4075;
    assign out10[51] = w4076;
    assign out10[52] = w4077;
    assign out10[53] = w4078;
    assign out10[54] = w4079;
    assign out10[55] = w4080;
    assign out10[56] = w4081;
    assign out10[57] = w4082;
    assign out10[58] = w4083;
    assign out10[59] = w4084;
    assign out10[60] = w4085;
    assign out10[61] = w4086;
    assign out10[62] = w4087;
    assign out10[63] = w4088;
    assign out10[64] = w4089;
    assign out10[65] = w4090;
    assign out10[66] = w4091;
    assign out10[67] = w4092;
    assign out10[68] = w4093;
    assign out10[69] = w4801;
    assign out10[70] = w4802;
    assign out10[71] = w4803;
    assign out10[72] = w4804;
    wire w2246;
    wire w2247;
    wire w2248;
    wire w2249;
    wire w2250;
    wire w2251;
    wire w2252;
    wire w2253;
    wire w2254;
    wire w2255;
    wire w2256;
    wire w2257;
    wire w2258;
    wire w2259;
    wire w2260;
    wire w2261;
    wire w2262;
    wire w2263;
    wire w2264;
    wire w2265;
    wire w2266;
    wire w2267;
    wire w2268;
    wire w2269;
    wire w2270;
    wire w2271;
    wire w2272;
    wire w2273;
    wire w2274;
    wire w2275;
    wire w2276;
    wire w2277;
    wire w2278;
    wire w2279;
    wire w2280;
    wire w2281;
    wire w2282;
    wire w2283;
    wire w2284;
    wire w2285;
    wire w2286;
    wire w2287;
    wire w2288;
    wire w2289;
    wire w2290;
    wire w2291;
    wire w2292;
    wire w2293;
    wire w2294;
    wire w2295;
    wire w2296;
    wire w2297;
    wire w2298;
    wire w2299;
    wire w2300;
    wire w2301;
    wire w2302;
    wire w2303;
    wire w2304;
    wire w2305;
    wire w2306;
    wire w2307;
    wire w2308;
    wire w2309;
    wire w2310;
    wire w2311;
    wire w2312;
    wire w2313;
    wire w2314;
    wire w4805;
    wire w4806;
    wire w4807;
    wire w4808;
    assign out11[0] = w2246;
    assign out11[1] = w2247;
    assign out11[2] = w2248;
    assign out11[3] = w2249;
    assign out11[4] = w2250;
    assign out11[5] = w2251;
    assign out11[6] = w2252;
    assign out11[7] = w2253;
    assign out11[8] = w2254;
    assign out11[9] = w2255;
    assign out11[10] = w2256;
    assign out11[11] = w2257;
    assign out11[12] = w2258;
    assign out11[13] = w2259;
    assign out11[14] = w2260;
    assign out11[15] = w2261;
    assign out11[16] = w2262;
    assign out11[17] = w2263;
    assign out11[18] = w2264;
    assign out11[19] = w2265;
    assign out11[20] = w2266;
    assign out11[21] = w2267;
    assign out11[22] = w2268;
    assign out11[23] = w2269;
    assign out11[24] = w2270;
    assign out11[25] = w2271;
    assign out11[26] = w2272;
    assign out11[27] = w2273;
    assign out11[28] = w2274;
    assign out11[29] = w2275;
    assign out11[30] = w2276;
    assign out11[31] = w2277;
    assign out11[32] = w2278;
    assign out11[33] = w2279;
    assign out11[34] = w2280;
    assign out11[35] = w2281;
    assign out11[36] = w2282;
    assign out11[37] = w2283;
    assign out11[38] = w2284;
    assign out11[39] = w2285;
    assign out11[40] = w2286;
    assign out11[41] = w2287;
    assign out11[42] = w2288;
    assign out11[43] = w2289;
    assign out11[44] = w2290;
    assign out11[45] = w2291;
    assign out11[46] = w2292;
    assign out11[47] = w2293;
    assign out11[48] = w2294;
    assign out11[49] = w2295;
    assign out11[50] = w2296;
    assign out11[51] = w2297;
    assign out11[52] = w2298;
    assign out11[53] = w2299;
    assign out11[54] = w2300;
    assign out11[55] = w2301;
    assign out11[56] = w2302;
    assign out11[57] = w2303;
    assign out11[58] = w2304;
    assign out11[59] = w2305;
    assign out11[60] = w2306;
    assign out11[61] = w2307;
    assign out11[62] = w2308;
    assign out11[63] = w2309;
    assign out11[64] = w2310;
    assign out11[65] = w2311;
    assign out11[66] = w2312;
    assign out11[67] = w2313;
    assign out11[68] = w2314;
    assign out11[69] = w4805;
    assign out11[70] = w4806;
    assign out11[71] = w4807;
    assign out11[72] = w4808;
    wire w4469;
    wire w4470;
    wire w4471;
    wire w4472;
    wire w4473;
    wire w4474;
    wire w4475;
    wire w4476;
    wire w4477;
    wire w4478;
    wire w4479;
    wire w4480;
    wire w4481;
    wire w4482;
    wire w4483;
    wire w4484;
    wire w4485;
    wire w4486;
    wire w4487;
    wire w4488;
    wire w4489;
    wire w4490;
    wire w4491;
    wire w4492;
    wire w4493;
    wire w4494;
    wire w4495;
    wire w4496;
    wire w4497;
    wire w4498;
    wire w4499;
    wire w4500;
    wire w4501;
    wire w4502;
    wire w4503;
    wire w4504;
    wire w4505;
    wire w4506;
    wire w4507;
    wire w4508;
    wire w4509;
    wire w4510;
    wire w4511;
    wire w4512;
    wire w4513;
    wire w4514;
    wire w4515;
    wire w4516;
    wire w4517;
    wire w4518;
    wire w4519;
    wire w4520;
    wire w4521;
    wire w4522;
    wire w4523;
    wire w4524;
    wire w4525;
    wire w4526;
    wire w4527;
    wire w4528;
    wire w4529;
    wire w4530;
    wire w4531;
    wire w4532;
    wire w4533;
    wire w4534;
    wire w4535;
    wire w4536;
    wire w4537;
    wire w4809;
    wire w4810;
    wire w4811;
    wire w4812;
    assign out12[0] = w4469;
    assign out12[1] = w4470;
    assign out12[2] = w4471;
    assign out12[3] = w4472;
    assign out12[4] = w4473;
    assign out12[5] = w4474;
    assign out12[6] = w4475;
    assign out12[7] = w4476;
    assign out12[8] = w4477;
    assign out12[9] = w4478;
    assign out12[10] = w4479;
    assign out12[11] = w4480;
    assign out12[12] = w4481;
    assign out12[13] = w4482;
    assign out12[14] = w4483;
    assign out12[15] = w4484;
    assign out12[16] = w4485;
    assign out12[17] = w4486;
    assign out12[18] = w4487;
    assign out12[19] = w4488;
    assign out12[20] = w4489;
    assign out12[21] = w4490;
    assign out12[22] = w4491;
    assign out12[23] = w4492;
    assign out12[24] = w4493;
    assign out12[25] = w4494;
    assign out12[26] = w4495;
    assign out12[27] = w4496;
    assign out12[28] = w4497;
    assign out12[29] = w4498;
    assign out12[30] = w4499;
    assign out12[31] = w4500;
    assign out12[32] = w4501;
    assign out12[33] = w4502;
    assign out12[34] = w4503;
    assign out12[35] = w4504;
    assign out12[36] = w4505;
    assign out12[37] = w4506;
    assign out12[38] = w4507;
    assign out12[39] = w4508;
    assign out12[40] = w4509;
    assign out12[41] = w4510;
    assign out12[42] = w4511;
    assign out12[43] = w4512;
    assign out12[44] = w4513;
    assign out12[45] = w4514;
    assign out12[46] = w4515;
    assign out12[47] = w4516;
    assign out12[48] = w4517;
    assign out12[49] = w4518;
    assign out12[50] = w4519;
    assign out12[51] = w4520;
    assign out12[52] = w4521;
    assign out12[53] = w4522;
    assign out12[54] = w4523;
    assign out12[55] = w4524;
    assign out12[56] = w4525;
    assign out12[57] = w4526;
    assign out12[58] = w4527;
    assign out12[59] = w4528;
    assign out12[60] = w4529;
    assign out12[61] = w4530;
    assign out12[62] = w4531;
    assign out12[63] = w4532;
    assign out12[64] = w4533;
    assign out12[65] = w4534;
    assign out12[66] = w4535;
    assign out12[67] = w4536;
    assign out12[68] = w4537;
    assign out12[69] = w4809;
    assign out12[70] = w4810;
    assign out12[71] = w4811;
    assign out12[72] = w4812;
    wire w2690;
    wire w2691;
    wire w2692;
    wire w2693;
    wire w2694;
    wire w2695;
    wire w2696;
    wire w2697;
    wire w2698;
    wire w2699;
    wire w2700;
    wire w2701;
    wire w2702;
    wire w2703;
    wire w2704;
    wire w2705;
    wire w2706;
    wire w2707;
    wire w2708;
    wire w2709;
    wire w2710;
    wire w2711;
    wire w2712;
    wire w2713;
    wire w2714;
    wire w2715;
    wire w2716;
    wire w2717;
    wire w2718;
    wire w2719;
    wire w2720;
    wire w2721;
    wire w2722;
    wire w2723;
    wire w2724;
    wire w2725;
    wire w2726;
    wire w2727;
    wire w2728;
    wire w2729;
    wire w2730;
    wire w2731;
    wire w2732;
    wire w2733;
    wire w2734;
    wire w2735;
    wire w2736;
    wire w2737;
    wire w2738;
    wire w2739;
    wire w2740;
    wire w2741;
    wire w2742;
    wire w2743;
    wire w2744;
    wire w2745;
    wire w2746;
    wire w2747;
    wire w2748;
    wire w2749;
    wire w2750;
    wire w2751;
    wire w2752;
    wire w2753;
    wire w2754;
    wire w2755;
    wire w2756;
    wire w2757;
    wire w2758;
    wire w4813;
    wire w4814;
    wire w4815;
    wire w4816;
    assign out13[0] = w2690;
    assign out13[1] = w2691;
    assign out13[2] = w2692;
    assign out13[3] = w2693;
    assign out13[4] = w2694;
    assign out13[5] = w2695;
    assign out13[6] = w2696;
    assign out13[7] = w2697;
    assign out13[8] = w2698;
    assign out13[9] = w2699;
    assign out13[10] = w2700;
    assign out13[11] = w2701;
    assign out13[12] = w2702;
    assign out13[13] = w2703;
    assign out13[14] = w2704;
    assign out13[15] = w2705;
    assign out13[16] = w2706;
    assign out13[17] = w2707;
    assign out13[18] = w2708;
    assign out13[19] = w2709;
    assign out13[20] = w2710;
    assign out13[21] = w2711;
    assign out13[22] = w2712;
    assign out13[23] = w2713;
    assign out13[24] = w2714;
    assign out13[25] = w2715;
    assign out13[26] = w2716;
    assign out13[27] = w2717;
    assign out13[28] = w2718;
    assign out13[29] = w2719;
    assign out13[30] = w2720;
    assign out13[31] = w2721;
    assign out13[32] = w2722;
    assign out13[33] = w2723;
    assign out13[34] = w2724;
    assign out13[35] = w2725;
    assign out13[36] = w2726;
    assign out13[37] = w2727;
    assign out13[38] = w2728;
    assign out13[39] = w2729;
    assign out13[40] = w2730;
    assign out13[41] = w2731;
    assign out13[42] = w2732;
    assign out13[43] = w2733;
    assign out13[44] = w2734;
    assign out13[45] = w2735;
    assign out13[46] = w2736;
    assign out13[47] = w2737;
    assign out13[48] = w2738;
    assign out13[49] = w2739;
    assign out13[50] = w2740;
    assign out13[51] = w2741;
    assign out13[52] = w2742;
    assign out13[53] = w2743;
    assign out13[54] = w2744;
    assign out13[55] = w2745;
    assign out13[56] = w2746;
    assign out13[57] = w2747;
    assign out13[58] = w2748;
    assign out13[59] = w2749;
    assign out13[60] = w2750;
    assign out13[61] = w2751;
    assign out13[62] = w2752;
    assign out13[63] = w2753;
    assign out13[64] = w2754;
    assign out13[65] = w2755;
    assign out13[66] = w2756;
    assign out13[67] = w2757;
    assign out13[68] = w2758;
    assign out13[69] = w4813;
    assign out13[70] = w4814;
    assign out13[71] = w4815;
    assign out13[72] = w4816;
    wire w3879;
    wire w3880;
    wire w3881;
    wire w3882;
    wire w3883;
    wire w3884;
    wire w3885;
    wire w3886;
    wire w3887;
    wire w3888;
    wire w3889;
    wire w3890;
    wire w3891;
    wire w3892;
    wire w3893;
    wire w3894;
    wire w3895;
    wire w3896;
    wire w3897;
    wire w3898;
    wire w3899;
    wire w3900;
    wire w3901;
    wire w3902;
    wire w3903;
    wire w3904;
    wire w3905;
    wire w3906;
    wire w3907;
    wire w3908;
    wire w3909;
    wire w3910;
    wire w3911;
    wire w3912;
    wire w3913;
    wire w3914;
    wire w3915;
    wire w3916;
    wire w3917;
    wire w3918;
    wire w3919;
    wire w3920;
    wire w3921;
    wire w3922;
    wire w3923;
    wire w3924;
    wire w3925;
    wire w3926;
    wire w3927;
    wire w3928;
    wire w3929;
    wire w3930;
    wire w3931;
    wire w3932;
    wire w3933;
    wire w3934;
    wire w3935;
    wire w3936;
    wire w3937;
    wire w3938;
    wire w3939;
    wire w3940;
    wire w3941;
    wire w3942;
    wire w3943;
    wire w3944;
    wire w3945;
    wire w3946;
    wire w3947;
    wire w4817;
    wire w4818;
    wire w4819;
    wire w4820;
    assign out14[0] = w3879;
    assign out14[1] = w3880;
    assign out14[2] = w3881;
    assign out14[3] = w3882;
    assign out14[4] = w3883;
    assign out14[5] = w3884;
    assign out14[6] = w3885;
    assign out14[7] = w3886;
    assign out14[8] = w3887;
    assign out14[9] = w3888;
    assign out14[10] = w3889;
    assign out14[11] = w3890;
    assign out14[12] = w3891;
    assign out14[13] = w3892;
    assign out14[14] = w3893;
    assign out14[15] = w3894;
    assign out14[16] = w3895;
    assign out14[17] = w3896;
    assign out14[18] = w3897;
    assign out14[19] = w3898;
    assign out14[20] = w3899;
    assign out14[21] = w3900;
    assign out14[22] = w3901;
    assign out14[23] = w3902;
    assign out14[24] = w3903;
    assign out14[25] = w3904;
    assign out14[26] = w3905;
    assign out14[27] = w3906;
    assign out14[28] = w3907;
    assign out14[29] = w3908;
    assign out14[30] = w3909;
    assign out14[31] = w3910;
    assign out14[32] = w3911;
    assign out14[33] = w3912;
    assign out14[34] = w3913;
    assign out14[35] = w3914;
    assign out14[36] = w3915;
    assign out14[37] = w3916;
    assign out14[38] = w3917;
    assign out14[39] = w3918;
    assign out14[40] = w3919;
    assign out14[41] = w3920;
    assign out14[42] = w3921;
    assign out14[43] = w3922;
    assign out14[44] = w3923;
    assign out14[45] = w3924;
    assign out14[46] = w3925;
    assign out14[47] = w3926;
    assign out14[48] = w3927;
    assign out14[49] = w3928;
    assign out14[50] = w3929;
    assign out14[51] = w3930;
    assign out14[52] = w3931;
    assign out14[53] = w3932;
    assign out14[54] = w3933;
    assign out14[55] = w3934;
    assign out14[56] = w3935;
    assign out14[57] = w3936;
    assign out14[58] = w3937;
    assign out14[59] = w3938;
    assign out14[60] = w3939;
    assign out14[61] = w3940;
    assign out14[62] = w3941;
    assign out14[63] = w3942;
    assign out14[64] = w3943;
    assign out14[65] = w3944;
    assign out14[66] = w3945;
    assign out14[67] = w3946;
    assign out14[68] = w3947;
    assign out14[69] = w4817;
    assign out14[70] = w4818;
    assign out14[71] = w4819;
    assign out14[72] = w4820;
    wire w2100;
    wire w2101;
    wire w2102;
    wire w2103;
    wire w2104;
    wire w2105;
    wire w2106;
    wire w2107;
    wire w2108;
    wire w2109;
    wire w2110;
    wire w2111;
    wire w2112;
    wire w2113;
    wire w2114;
    wire w2115;
    wire w2116;
    wire w2117;
    wire w2118;
    wire w2119;
    wire w2120;
    wire w2121;
    wire w2122;
    wire w2123;
    wire w2124;
    wire w2125;
    wire w2126;
    wire w2127;
    wire w2128;
    wire w2129;
    wire w2130;
    wire w2131;
    wire w2132;
    wire w2133;
    wire w2134;
    wire w2135;
    wire w2136;
    wire w2137;
    wire w2138;
    wire w2139;
    wire w2140;
    wire w2141;
    wire w2142;
    wire w2143;
    wire w2144;
    wire w2145;
    wire w2146;
    wire w2147;
    wire w2148;
    wire w2149;
    wire w2150;
    wire w2151;
    wire w2152;
    wire w2153;
    wire w2154;
    wire w2155;
    wire w2156;
    wire w2157;
    wire w2158;
    wire w2159;
    wire w2160;
    wire w2161;
    wire w2162;
    wire w2163;
    wire w2164;
    wire w2165;
    wire w2166;
    wire w2167;
    wire w2168;
    wire w4821;
    wire w4822;
    wire w4823;
    wire w4824;
    assign out15[0] = w2100;
    assign out15[1] = w2101;
    assign out15[2] = w2102;
    assign out15[3] = w2103;
    assign out15[4] = w2104;
    assign out15[5] = w2105;
    assign out15[6] = w2106;
    assign out15[7] = w2107;
    assign out15[8] = w2108;
    assign out15[9] = w2109;
    assign out15[10] = w2110;
    assign out15[11] = w2111;
    assign out15[12] = w2112;
    assign out15[13] = w2113;
    assign out15[14] = w2114;
    assign out15[15] = w2115;
    assign out15[16] = w2116;
    assign out15[17] = w2117;
    assign out15[18] = w2118;
    assign out15[19] = w2119;
    assign out15[20] = w2120;
    assign out15[21] = w2121;
    assign out15[22] = w2122;
    assign out15[23] = w2123;
    assign out15[24] = w2124;
    assign out15[25] = w2125;
    assign out15[26] = w2126;
    assign out15[27] = w2127;
    assign out15[28] = w2128;
    assign out15[29] = w2129;
    assign out15[30] = w2130;
    assign out15[31] = w2131;
    assign out15[32] = w2132;
    assign out15[33] = w2133;
    assign out15[34] = w2134;
    assign out15[35] = w2135;
    assign out15[36] = w2136;
    assign out15[37] = w2137;
    assign out15[38] = w2138;
    assign out15[39] = w2139;
    assign out15[40] = w2140;
    assign out15[41] = w2141;
    assign out15[42] = w2142;
    assign out15[43] = w2143;
    assign out15[44] = w2144;
    assign out15[45] = w2145;
    assign out15[46] = w2146;
    assign out15[47] = w2147;
    assign out15[48] = w2148;
    assign out15[49] = w2149;
    assign out15[50] = w2150;
    assign out15[51] = w2151;
    assign out15[52] = w2152;
    assign out15[53] = w2153;
    assign out15[54] = w2154;
    assign out15[55] = w2155;
    assign out15[56] = w2156;
    assign out15[57] = w2157;
    assign out15[58] = w2158;
    assign out15[59] = w2159;
    assign out15[60] = w2160;
    assign out15[61] = w2161;
    assign out15[62] = w2162;
    assign out15[63] = w2163;
    assign out15[64] = w2164;
    assign out15[65] = w2165;
    assign out15[66] = w2166;
    assign out15[67] = w2167;
    assign out15[68] = w2168;
    assign out15[69] = w4821;
    assign out15[70] = w4822;
    assign out15[71] = w4823;
    assign out15[72] = w4824;
    wire w6;
    xor xor0(w6, x11_68, x12_68);
    wire w7;
    xor xor1(w7, x13_68, x14_68);
    wire w1;
    xor xor2(w1, x1_68, x2_68);
    wire w2;
    xor xor3(w2, x3_68, x4_68);
    wire w3;
    xor xor4(w3, x5_68, x6_68);
    wire w4;
    xor xor5(w4, x7_68, x8_68);
    wire w5;
    xor xor6(w5, x9_68, x10_68);
    wire w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99;
    sw_m #(.SIZE(74)) sw7({w92,w91,w90,w89,w88,w87,w86,w85,w84,w83,w82,w81,w80,w79,w78,w77,w76,w75,w74,w73,w72,w71,w70,w69,w68,w67,w66,w65,w64,w63,w62,w61,w60,w59,w58,w57,w56,w55,w54,w53,w52,w51,w50,w49,w48,w47,w46,w45,w44,w43,w42,w41,w40,w39,w38,w37,w36,w35,w34,w33,w32,w31,w30,w29,w28,w27,w26,w25,w24,w23,w22,w21,w20,w19}, {w166,w165,w164,w163,w162,w161,w160,w159,w158,w157,w156,w155,w154,w153,w152,w151,w150,w149,w148,w147,w146,w145,w144,w143,w142,w141,w140,w139,w138,w137,w136,w135,w134,w133,w132,w131,w130,w129,w128,w127,w126,w125,w124,w123,w122,w121,w120,w119,w118,w117,w116,w115,w114,w113,w112,w111,w110,w109,w108,w107,w106,w105,w104,w103,w102,w101,w100,w99,w98,w97,w96,w95,w94,w93}, x0_68, {x0_68,x0_72,x0_71,x0_70,x0_69,x0_68,x0_67,x0_66,x0_65,x0_64,x0_63,x0_62,x0_61,x0_60,x0_59,x0_58,x0_57,x0_56,x0_55,x0_54,x0_53,x0_52,x0_51,x0_50,x0_49,x0_48,x0_47,x0_46,x0_45,x0_44,x0_43,x0_42,x0_41,x0_40,x0_39,x0_38,x0_37,x0_36,x0_35,x0_34,x0_33,x0_32,x0_31,x0_30,x0_29,x0_28,x0_27,x0_26,x0_25,x0_24,x0_23,x0_22,x0_21,x0_20,x0_19,x0_18,x0_17,x0_16,x0_15,x0_14,x0_13,x0_12,x0_11,x0_10,x0_9,x0_8,x0_7,x0_6,x0_5,x0_4,x0_3,x0_2,x0_1,x0_0}, {x1_68,x1_72,x1_71,x1_70,x1_69,x1_68,x1_67,x1_66,x1_65,x1_64,x1_63,x1_62,x1_61,x1_60,x1_59,x1_58,x1_57,x1_56,x1_55,x1_54,x1_53,x1_52,x1_51,x1_50,x1_49,x1_48,x1_47,x1_46,x1_45,x1_44,x1_43,x1_42,x1_41,x1_40,x1_39,x1_38,x1_37,x1_36,x1_35,x1_34,x1_33,x1_32,x1_31,x1_30,x1_29,x1_28,x1_27,x1_26,x1_25,x1_24,x1_23,x1_22,x1_21,x1_20,x1_19,x1_18,x1_17,x1_16,x1_15,x1_14,x1_13,x1_12,x1_11,x1_10,x1_9,x1_8,x1_7,x1_6,x1_5,x1_4,x1_3,x1_2,x1_1,x1_0});
    wire w9;
    xor xor8(w9, w2, w3);
    wire w10;
    xor xor9(w10, w4, w5);
    wire w11;
    xor xor10(w11, w6, w7);
    wire w8;
    xor xor11(w8, x0_68, w1);
    wire w13;
    xor xor12(w13, w10, w11);
    wire w16;
    xor xor13(w16, w8, w2);
    wire w12;
    xor xor14(w12, w8, w9);
    wire w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314;
    sw_m #(.SIZE(74)) sw15({w240,w239,w238,w237,w236,w235,w234,w233,w232,w231,w230,w229,w228,w227,w226,w225,w224,w223,w222,w221,w220,w219,w218,w217,w216,w215,w214,w213,w212,w211,w210,w209,w208,w207,w206,w205,w204,w203,w202,w201,w200,w199,w198,w197,w196,w195,w194,w193,w192,w191,w190,w189,w188,w187,w186,w185,w184,w183,w182,w181,w180,w179,w178,w177,w176,w175,w174,w173,w172,w171,w170,w169,w168,w167}, {w314,w313,w312,w311,w310,w309,w308,w307,w306,w305,w304,w303,w302,w301,w300,w299,w298,w297,w296,w295,w294,w293,w292,w291,w290,w289,w288,w287,w286,w285,w284,w283,w282,w281,w280,w279,w278,w277,w276,w275,w274,w273,w272,w271,w270,w269,w268,w267,w266,w265,w264,w263,w262,w261,w260,w259,w258,w257,w256,w255,w254,w253,w252,w251,w250,w249,w248,w247,w246,w245,w244,w243,w242,w241}, w8, {x2_68,x2_72,x2_71,x2_70,x2_69,x2_68,x2_67,x2_66,x2_65,x2_64,x2_63,x2_62,x2_61,x2_60,x2_59,x2_58,x2_57,x2_56,x2_55,x2_54,x2_53,x2_52,x2_51,x2_50,x2_49,x2_48,x2_47,x2_46,x2_45,x2_44,x2_43,x2_42,x2_41,x2_40,x2_39,x2_38,x2_37,x2_36,x2_35,x2_34,x2_33,x2_32,x2_31,x2_30,x2_29,x2_28,x2_27,x2_26,x2_25,x2_24,x2_23,x2_22,x2_21,x2_20,x2_19,x2_18,x2_17,x2_16,x2_15,x2_14,x2_13,x2_12,x2_11,x2_10,x2_9,x2_8,x2_7,x2_6,x2_5,x2_4,x2_3,x2_2,x2_1,x2_0}, {x3_68,x3_72,x3_71,x3_70,x3_69,x3_68,x3_67,x3_66,x3_65,x3_64,x3_63,x3_62,x3_61,x3_60,x3_59,x3_58,x3_57,x3_56,x3_55,x3_54,x3_53,x3_52,x3_51,x3_50,x3_49,x3_48,x3_47,x3_46,x3_45,x3_44,x3_43,x3_42,x3_41,x3_40,x3_39,x3_38,x3_37,x3_36,x3_35,x3_34,x3_33,x3_32,x3_31,x3_30,x3_29,x3_28,x3_27,x3_26,x3_25,x3_24,x3_23,x3_22,x3_21,x3_20,x3_19,x3_18,x3_17,x3_16,x3_15,x3_14,x3_13,x3_12,x3_11,x3_10,x3_9,x3_8,x3_7,x3_6,x3_5,x3_4,x3_3,x3_2,x3_1,x3_0});
    wire w15;
    xor xor16(w15, w12, w10);
    wire w14;
    xor xor17(w14, w12, w13);
    wire w17;
    xor xor18(w17, w12, w4);
    wire w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610;
    sw_m #(.SIZE(74)) sw19({w536,w535,w534,w533,w532,w531,w530,w529,w528,w527,w526,w525,w524,w523,w522,w521,w520,w519,w518,w517,w516,w515,w514,w513,w512,w511,w510,w509,w508,w507,w506,w505,w504,w503,w502,w501,w500,w499,w498,w497,w496,w495,w494,w493,w492,w491,w490,w489,w488,w487,w486,w485,w484,w483,w482,w481,w480,w479,w478,w477,w476,w475,w474,w473,w472,w471,w470,w469,w468,w467,w466,w465,w464,w463}, {w610,w609,w608,w607,w606,w605,w604,w603,w602,w601,w600,w599,w598,w597,w596,w595,w594,w593,w592,w591,w590,w589,w588,w587,w586,w585,w584,w583,w582,w581,w580,w579,w578,w577,w576,w575,w574,w573,w572,w571,w570,w569,w568,w567,w566,w565,w564,w563,w562,w561,w560,w559,w558,w557,w556,w555,w554,w553,w552,w551,w550,w549,w548,w547,w546,w545,w544,w543,w542,w541,w540,w539,w538,w537}, w12, {x6_68,x6_72,x6_71,x6_70,x6_69,x6_68,x6_67,x6_66,x6_65,x6_64,x6_63,x6_62,x6_61,x6_60,x6_59,x6_58,x6_57,x6_56,x6_55,x6_54,x6_53,x6_52,x6_51,x6_50,x6_49,x6_48,x6_47,x6_46,x6_45,x6_44,x6_43,x6_42,x6_41,x6_40,x6_39,x6_38,x6_37,x6_36,x6_35,x6_34,x6_33,x6_32,x6_31,x6_30,x6_29,x6_28,x6_27,x6_26,x6_25,x6_24,x6_23,x6_22,x6_21,x6_20,x6_19,x6_18,x6_17,x6_16,x6_15,x6_14,x6_13,x6_12,x6_11,x6_10,x6_9,x6_8,x6_7,x6_6,x6_5,x6_4,x6_3,x6_2,x6_1,x6_0}, {x7_68,x7_72,x7_71,x7_70,x7_69,x7_68,x7_67,x7_66,x7_65,x7_64,x7_63,x7_62,x7_61,x7_60,x7_59,x7_58,x7_57,x7_56,x7_55,x7_54,x7_53,x7_52,x7_51,x7_50,x7_49,x7_48,x7_47,x7_46,x7_45,x7_44,x7_43,x7_42,x7_41,x7_40,x7_39,x7_38,x7_37,x7_36,x7_35,x7_34,x7_33,x7_32,x7_31,x7_30,x7_29,x7_28,x7_27,x7_26,x7_25,x7_24,x7_23,x7_22,x7_21,x7_20,x7_19,x7_18,x7_17,x7_16,x7_15,x7_14,x7_13,x7_12,x7_11,x7_10,x7_9,x7_8,x7_7,x7_6,x7_5,x7_4,x7_3,x7_2,x7_1,x7_0});
    wire w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462;
    sw_m #(.SIZE(74)) sw20({w388,w387,w386,w385,w384,w383,w382,w381,w380,w379,w378,w377,w376,w375,w374,w373,w372,w371,w370,w369,w368,w367,w366,w365,w364,w363,w362,w361,w360,w359,w358,w357,w356,w355,w354,w353,w352,w351,w350,w349,w348,w347,w346,w345,w344,w343,w342,w341,w340,w339,w338,w337,w336,w335,w334,w333,w332,w331,w330,w329,w328,w327,w326,w325,w324,w323,w322,w321,w320,w319,w318,w317,w316,w315}, {w462,w461,w460,w459,w458,w457,w456,w455,w454,w453,w452,w451,w450,w449,w448,w447,w446,w445,w444,w443,w442,w441,w440,w439,w438,w437,w436,w435,w434,w433,w432,w431,w430,w429,w428,w427,w426,w425,w424,w423,w422,w421,w420,w419,w418,w417,w416,w415,w414,w413,w412,w411,w410,w409,w408,w407,w406,w405,w404,w403,w402,w401,w400,w399,w398,w397,w396,w395,w394,w393,w392,w391,w390,w389}, w16, {x4_68,x4_72,x4_71,x4_70,x4_69,x4_68,x4_67,x4_66,x4_65,x4_64,x4_63,x4_62,x4_61,x4_60,x4_59,x4_58,x4_57,x4_56,x4_55,x4_54,x4_53,x4_52,x4_51,x4_50,x4_49,x4_48,x4_47,x4_46,x4_45,x4_44,x4_43,x4_42,x4_41,x4_40,x4_39,x4_38,x4_37,x4_36,x4_35,x4_34,x4_33,x4_32,x4_31,x4_30,x4_29,x4_28,x4_27,x4_26,x4_25,x4_24,x4_23,x4_22,x4_21,x4_20,x4_19,x4_18,x4_17,x4_16,x4_15,x4_14,x4_13,x4_12,x4_11,x4_10,x4_9,x4_8,x4_7,x4_6,x4_5,x4_4,x4_3,x4_2,x4_1,x4_0}, {x5_68,x5_72,x5_71,x5_70,x5_69,x5_68,x5_67,x5_66,x5_65,x5_64,x5_63,x5_62,x5_61,x5_60,x5_59,x5_58,x5_57,x5_56,x5_55,x5_54,x5_53,x5_52,x5_51,x5_50,x5_49,x5_48,x5_47,x5_46,x5_45,x5_44,x5_43,x5_42,x5_41,x5_40,x5_39,x5_38,x5_37,x5_36,x5_35,x5_34,x5_33,x5_32,x5_31,x5_30,x5_29,x5_28,x5_27,x5_26,x5_25,x5_24,x5_23,x5_22,x5_21,x5_20,x5_19,x5_18,x5_17,x5_16,x5_15,x5_14,x5_13,x5_12,x5_11,x5_10,x5_9,x5_8,x5_7,x5_6,x5_5,x5_4,x5_3,x5_2,x5_1,x5_0});
    wire w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136;
    sw_m #(.SIZE(74)) sw21({w3062,w3061,w3060,w3059,w3058,w3057,w3056,w3055,w3054,w3053,w3052,w3051,w3050,w3049,w3048,w3047,w3046,w3045,w3044,w3043,w3042,w3041,w3040,w3039,w3038,w3037,w3036,w3035,w3034,w3033,w3032,w3031,w3030,w3029,w3028,w3027,w3026,w3025,w3024,w3023,w3022,w3021,w3020,w3019,w3018,w3017,w3016,w3015,w3014,w3013,w3012,w3011,w3010,w3009,w3008,w3007,w3006,w3005,w3004,w3003,w3002,w3001,w3000,w2999,w2998,w2997,w2996,w2995,w2994,w2993,w2992,w2991,w2990,w2989}, {w3136,w3135,w3134,w3133,w3132,w3131,w3130,w3129,w3128,w3127,w3126,w3125,w3124,w3123,w3122,w3121,w3120,w3119,w3118,w3117,w3116,w3115,w3114,w3113,w3112,w3111,w3110,w3109,w3108,w3107,w3106,w3105,w3104,w3103,w3102,w3101,w3100,w3099,w3098,w3097,w3096,w3095,w3094,w3093,w3092,w3091,w3090,w3089,w3088,w3087,w3086,w3085,w3084,w3083,w3082,w3081,w3080,w3079,w3078,w3077,w3076,w3075,w3074,w3073,w3072,w3071,w3070,w3069,w3068,w3067,w3066,w3065,w3064,w3063}, w166, {w166,w165,w164,w163,w162,w161,w160,w159,w158,w157,w156,w155,w154,w153,w152,w151,w150,w149,w148,w147,w146,w145,w144,w143,w142,w141,w140,w139,w138,w137,w136,w135,w134,w133,w132,w131,w130,w129,w128,w127,w126,w125,w124,w123,w122,w121,w120,w119,w118,w117,w116,w115,w114,w113,w112,w111,w110,w109,w108,w107,w106,w105,w104,w103,w102,w101,w100,w99,w98,w97,w96,w95,w94,w93}, {w314,w313,w312,w311,w310,w309,w308,w307,w306,w305,w304,w303,w302,w301,w300,w299,w298,w297,w296,w295,w294,w293,w292,w291,w290,w289,w288,w287,w286,w285,w284,w283,w282,w281,w280,w279,w278,w277,w276,w275,w274,w273,w272,w271,w270,w269,w268,w267,w266,w265,w264,w263,w262,w261,w260,w259,w258,w257,w256,w255,w254,w253,w252,w251,w250,w249,w248,w247,w246,w245,w244,w243,w242,w241});
    wire w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357;
    sw_m #(.SIZE(74)) sw22({w1283,w1282,w1281,w1280,w1279,w1278,w1277,w1276,w1275,w1274,w1273,w1272,w1271,w1270,w1269,w1268,w1267,w1266,w1265,w1264,w1263,w1262,w1261,w1260,w1259,w1258,w1257,w1256,w1255,w1254,w1253,w1252,w1251,w1250,w1249,w1248,w1247,w1246,w1245,w1244,w1243,w1242,w1241,w1240,w1239,w1238,w1237,w1236,w1235,w1234,w1233,w1232,w1231,w1230,w1229,w1228,w1227,w1226,w1225,w1224,w1223,w1222,w1221,w1220,w1219,w1218,w1217,w1216,w1215,w1214,w1213,w1212,w1211,w1210}, {w1357,w1356,w1355,w1354,w1353,w1352,w1351,w1350,w1349,w1348,w1347,w1346,w1345,w1344,w1343,w1342,w1341,w1340,w1339,w1338,w1337,w1336,w1335,w1334,w1333,w1332,w1331,w1330,w1329,w1328,w1327,w1326,w1325,w1324,w1323,w1322,w1321,w1320,w1319,w1318,w1317,w1316,w1315,w1314,w1313,w1312,w1311,w1310,w1309,w1308,w1307,w1306,w1305,w1304,w1303,w1302,w1301,w1300,w1299,w1298,w1297,w1296,w1295,w1294,w1293,w1292,w1291,w1290,w1289,w1288,w1287,w1286,w1285,w1284}, w92, {w92,w91,w90,w89,w88,w87,w86,w85,w84,w83,w82,w81,w80,w79,w78,w77,w76,w75,w74,w73,w72,w71,w70,w69,w68,w67,w66,w65,w64,w63,w62,w61,w60,w59,w58,w57,w56,w55,w54,w53,w52,w51,w50,w49,w48,w47,w46,w45,w44,w43,w42,w41,w40,w39,w38,w37,w36,w35,w34,w33,w32,w31,w30,w29,w28,w27,w26,w25,w24,w23,w22,w21,w20,w19}, {w240,w239,w238,w237,w236,w235,w234,w233,w232,w231,w230,w229,w228,w227,w226,w225,w224,w223,w222,w221,w220,w219,w218,w217,w216,w215,w214,w213,w212,w211,w210,w209,w208,w207,w206,w205,w204,w203,w202,w201,w200,w199,w198,w197,w196,w195,w194,w193,w192,w191,w190,w189,w188,w187,w186,w185,w184,w183,w182,w181,w180,w179,w178,w177,w176,w175,w174,w173,w172,w171,w170,w169,w168,w167});
    wire w18;
    xor xor23(w18, w15, w6);
    wire w1203;
    xor xor24(w1203, w240, w388);
    wire w2982;
    xor xor25(w2982, w314, w462);
    wire w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202;
    sw_m #(.SIZE(74)) sw26({w1128,w1127,w1126,w1125,w1124,w1123,w1122,w1121,w1120,w1119,w1118,w1117,w1116,w1115,w1114,w1113,w1112,w1111,w1110,w1109,w1108,w1107,w1106,w1105,w1104,w1103,w1102,w1101,w1100,w1099,w1098,w1097,w1096,w1095,w1094,w1093,w1092,w1091,w1090,w1089,w1088,w1087,w1086,w1085,w1084,w1083,w1082,w1081,w1080,w1079,w1078,w1077,w1076,w1075,w1074,w1073,w1072,w1071,w1070,w1069,w1068,w1067,w1066,w1065,w1064,w1063,w1062,w1061,w1060,w1059,w1058,w1057,w1056,w1055}, {w1202,w1201,w1200,w1199,w1198,w1197,w1196,w1195,w1194,w1193,w1192,w1191,w1190,w1189,w1188,w1187,w1186,w1185,w1184,w1183,w1182,w1181,w1180,w1179,w1178,w1177,w1176,w1175,w1174,w1173,w1172,w1171,w1170,w1169,w1168,w1167,w1166,w1165,w1164,w1163,w1162,w1161,w1160,w1159,w1158,w1157,w1156,w1155,w1154,w1153,w1152,w1151,w1150,w1149,w1148,w1147,w1146,w1145,w1144,w1143,w1142,w1141,w1140,w1139,w1138,w1137,w1136,w1135,w1134,w1133,w1132,w1131,w1130,w1129}, w14, {x14_68,x14_72,x14_71,x14_70,x14_69,x14_68,x14_67,x14_66,x14_65,x14_64,x14_63,x14_62,x14_61,x14_60,x14_59,x14_58,x14_57,x14_56,x14_55,x14_54,x14_53,x14_52,x14_51,x14_50,x14_49,x14_48,x14_47,x14_46,x14_45,x14_44,x14_43,x14_42,x14_41,x14_40,x14_39,x14_38,x14_37,x14_36,x14_35,x14_34,x14_33,x14_32,x14_31,x14_30,x14_29,x14_28,x14_27,x14_26,x14_25,x14_24,x14_23,x14_22,x14_21,x14_20,x14_19,x14_18,x14_17,x14_16,x14_15,x14_14,x14_13,x14_12,x14_11,x14_10,x14_9,x14_8,x14_7,x14_6,x14_5,x14_4,x14_3,x14_2,x14_1,x14_0}, {x15_68,x15_72,x15_71,x15_70,x15_69,x15_68,x15_67,x15_66,x15_65,x15_64,x15_63,x15_62,x15_61,x15_60,x15_59,x15_58,x15_57,x15_56,x15_55,x15_54,x15_53,x15_52,x15_51,x15_50,x15_49,x15_48,x15_47,x15_46,x15_45,x15_44,x15_43,x15_42,x15_41,x15_40,x15_39,x15_38,x15_37,x15_36,x15_35,x15_34,x15_33,x15_32,x15_31,x15_30,x15_29,x15_28,x15_27,x15_26,x15_25,x15_24,x15_23,x15_22,x15_21,x15_20,x15_19,x15_18,x15_17,x15_16,x15_15,x15_14,x15_13,x15_12,x15_11,x15_10,x15_9,x15_8,x15_7,x15_6,x15_5,x15_4,x15_3,x15_2,x15_1,x15_0});
    wire w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906;
    sw_m #(.SIZE(74)) sw27({w832,w831,w830,w829,w828,w827,w826,w825,w824,w823,w822,w821,w820,w819,w818,w817,w816,w815,w814,w813,w812,w811,w810,w809,w808,w807,w806,w805,w804,w803,w802,w801,w800,w799,w798,w797,w796,w795,w794,w793,w792,w791,w790,w789,w788,w787,w786,w785,w784,w783,w782,w781,w780,w779,w778,w777,w776,w775,w774,w773,w772,w771,w770,w769,w768,w767,w766,w765,w764,w763,w762,w761,w760,w759}, {w906,w905,w904,w903,w902,w901,w900,w899,w898,w897,w896,w895,w894,w893,w892,w891,w890,w889,w888,w887,w886,w885,w884,w883,w882,w881,w880,w879,w878,w877,w876,w875,w874,w873,w872,w871,w870,w869,w868,w867,w866,w865,w864,w863,w862,w861,w860,w859,w858,w857,w856,w855,w854,w853,w852,w851,w850,w849,w848,w847,w846,w845,w844,w843,w842,w841,w840,w839,w838,w837,w836,w835,w834,w833}, w15, {x10_68,x10_72,x10_71,x10_70,x10_69,x10_68,x10_67,x10_66,x10_65,x10_64,x10_63,x10_62,x10_61,x10_60,x10_59,x10_58,x10_57,x10_56,x10_55,x10_54,x10_53,x10_52,x10_51,x10_50,x10_49,x10_48,x10_47,x10_46,x10_45,x10_44,x10_43,x10_42,x10_41,x10_40,x10_39,x10_38,x10_37,x10_36,x10_35,x10_34,x10_33,x10_32,x10_31,x10_30,x10_29,x10_28,x10_27,x10_26,x10_25,x10_24,x10_23,x10_22,x10_21,x10_20,x10_19,x10_18,x10_17,x10_16,x10_15,x10_14,x10_13,x10_12,x10_11,x10_10,x10_9,x10_8,x10_7,x10_6,x10_5,x10_4,x10_3,x10_2,x10_1,x10_0}, {x11_68,x11_72,x11_71,x11_70,x11_69,x11_68,x11_67,x11_66,x11_65,x11_64,x11_63,x11_62,x11_61,x11_60,x11_59,x11_58,x11_57,x11_56,x11_55,x11_54,x11_53,x11_52,x11_51,x11_50,x11_49,x11_48,x11_47,x11_46,x11_45,x11_44,x11_43,x11_42,x11_41,x11_40,x11_39,x11_38,x11_37,x11_36,x11_35,x11_34,x11_33,x11_32,x11_31,x11_30,x11_29,x11_28,x11_27,x11_26,x11_25,x11_24,x11_23,x11_22,x11_21,x11_20,x11_19,x11_18,x11_17,x11_16,x11_15,x11_14,x11_13,x11_12,x11_11,x11_10,x11_9,x11_8,x11_7,x11_6,x11_5,x11_4,x11_3,x11_2,x11_1,x11_0});
    wire w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758;
    sw_m #(.SIZE(74)) sw28({w684,w683,w682,w681,w680,w679,w678,w677,w676,w675,w674,w673,w672,w671,w670,w669,w668,w667,w666,w665,w664,w663,w662,w661,w660,w659,w658,w657,w656,w655,w654,w653,w652,w651,w650,w649,w648,w647,w646,w645,w644,w643,w642,w641,w640,w639,w638,w637,w636,w635,w634,w633,w632,w631,w630,w629,w628,w627,w626,w625,w624,w623,w622,w621,w620,w619,w618,w617,w616,w615,w614,w613,w612,w611}, {w758,w757,w756,w755,w754,w753,w752,w751,w750,w749,w748,w747,w746,w745,w744,w743,w742,w741,w740,w739,w738,w737,w736,w735,w734,w733,w732,w731,w730,w729,w728,w727,w726,w725,w724,w723,w722,w721,w720,w719,w718,w717,w716,w715,w714,w713,w712,w711,w710,w709,w708,w707,w706,w705,w704,w703,w702,w701,w700,w699,w698,w697,w696,w695,w694,w693,w692,w691,w690,w689,w688,w687,w686,w685}, w17, {x8_68,x8_72,x8_71,x8_70,x8_69,x8_68,x8_67,x8_66,x8_65,x8_64,x8_63,x8_62,x8_61,x8_60,x8_59,x8_58,x8_57,x8_56,x8_55,x8_54,x8_53,x8_52,x8_51,x8_50,x8_49,x8_48,x8_47,x8_46,x8_45,x8_44,x8_43,x8_42,x8_41,x8_40,x8_39,x8_38,x8_37,x8_36,x8_35,x8_34,x8_33,x8_32,x8_31,x8_30,x8_29,x8_28,x8_27,x8_26,x8_25,x8_24,x8_23,x8_22,x8_21,x8_20,x8_19,x8_18,x8_17,x8_16,x8_15,x8_14,x8_13,x8_12,x8_11,x8_10,x8_9,x8_8,x8_7,x8_6,x8_5,x8_4,x8_3,x8_2,x8_1,x8_0}, {x9_68,x9_72,x9_71,x9_70,x9_69,x9_68,x9_67,x9_66,x9_65,x9_64,x9_63,x9_62,x9_61,x9_60,x9_59,x9_58,x9_57,x9_56,x9_55,x9_54,x9_53,x9_52,x9_51,x9_50,x9_49,x9_48,x9_47,x9_46,x9_45,x9_44,x9_43,x9_42,x9_41,x9_40,x9_39,x9_38,x9_37,x9_36,x9_35,x9_34,x9_33,x9_32,x9_31,x9_30,x9_29,x9_28,x9_27,x9_26,x9_25,x9_24,x9_23,x9_22,x9_21,x9_20,x9_19,x9_18,x9_17,x9_16,x9_15,x9_14,x9_13,x9_12,x9_11,x9_10,x9_9,x9_8,x9_7,x9_6,x9_5,x9_4,x9_3,x9_2,x9_1,x9_0});
    wire w2985;
    xor xor29(w2985, w166, w2982);
    wire w1204;
    xor xor30(w1204, w536, w684);
    wire w2983;
    xor xor31(w2983, w610, w758);
    wire w1206;
    xor xor32(w1206, w92, w1203);
    wire w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999;
    sw_m #(.SIZE(74)) sw33({w980,w979,w978,w977,w976,w975,w974,w973,w972,w971,w970,w969,w968,w967,w966,w965,w964,w963,w962,w961,w960,w959,w958,w957,w956,w955,w954,w953,w952,w951,w950,w949,w948,w947,w946,w945,w944,w943,w942,w941,w940,w939,w938,w937,w936,w935,w934,w933,w932,w931,w930,w929,w928,w927,w926,w925,w924,w923,w922,w921,w920,w919,w918,w917,w916,w915,w914,w913,w912,w911,w910,w909,w908,w907}, {w1054,w1053,w1052,w1051,w1050,w1049,w1048,w1047,w1046,w1045,w1044,w1043,w1042,w1041,w1040,w1039,w1038,w1037,w1036,w1035,w1034,w1033,w1032,w1031,w1030,w1029,w1028,w1027,w1026,w1025,w1024,w1023,w1022,w1021,w1020,w1019,w1018,w1017,w1016,w1015,w1014,w1013,w1012,w1011,w1010,w1009,w1008,w1007,w1006,w1005,w1004,w1003,w1002,w1001,w1000,w999,w998,w997,w996,w995,w994,w993,w992,w991,w990,w989,w988,w987,w986,w985,w984,w983,w982,w981}, w18, {x12_68,x12_72,x12_71,x12_70,x12_69,x12_68,x12_67,x12_66,x12_65,x12_64,x12_63,x12_62,x12_61,x12_60,x12_59,x12_58,x12_57,x12_56,x12_55,x12_54,x12_53,x12_52,x12_51,x12_50,x12_49,x12_48,x12_47,x12_46,x12_45,x12_44,x12_43,x12_42,x12_41,x12_40,x12_39,x12_38,x12_37,x12_36,x12_35,x12_34,x12_33,x12_32,x12_31,x12_30,x12_29,x12_28,x12_27,x12_26,x12_25,x12_24,x12_23,x12_22,x12_21,x12_20,x12_19,x12_18,x12_17,x12_16,x12_15,x12_14,x12_13,x12_12,x12_11,x12_10,x12_9,x12_8,x12_7,x12_6,x12_5,x12_4,x12_3,x12_2,x12_1,x12_0}, {x13_68,x13_72,x13_71,x13_70,x13_69,x13_68,x13_67,x13_66,x13_65,x13_64,x13_63,x13_62,x13_61,x13_60,x13_59,x13_58,x13_57,x13_56,x13_55,x13_54,x13_53,x13_52,x13_51,x13_50,x13_49,x13_48,x13_47,x13_46,x13_45,x13_44,x13_43,x13_42,x13_41,x13_40,x13_39,x13_38,x13_37,x13_36,x13_35,x13_34,x13_33,x13_32,x13_31,x13_30,x13_29,x13_28,x13_27,x13_26,x13_25,x13_24,x13_23,x13_22,x13_21,x13_20,x13_19,x13_18,x13_17,x13_16,x13_15,x13_14,x13_13,x13_12,x13_11,x13_10,x13_9,x13_8,x13_7,x13_6,x13_5,x13_4,x13_3,x13_2,x13_1,x13_0});
    wire w1209;
    xor xor34(w1209, w1206, w1204);
    wire w2988;
    xor xor35(w2988, w2985, w2983);
    wire w1205;
    xor xor36(w1205, w832, w980);
    wire w2984;
    xor xor37(w2984, w906, w1054);
    wire w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505;
    sw_m #(.SIZE(74)) sw38({w1431,w1430,w1429,w1428,w1427,w1426,w1425,w1424,w1423,w1422,w1421,w1420,w1419,w1418,w1417,w1416,w1415,w1414,w1413,w1412,w1411,w1410,w1409,w1408,w1407,w1406,w1405,w1404,w1403,w1402,w1401,w1400,w1399,w1398,w1397,w1396,w1395,w1394,w1393,w1392,w1391,w1390,w1389,w1388,w1387,w1386,w1385,w1384,w1383,w1382,w1381,w1380,w1379,w1378,w1377,w1376,w1375,w1374,w1373,w1372,w1371,w1370,w1369,w1368,w1367,w1366,w1365,w1364,w1363,w1362,w1361,w1360,w1359,w1358}, {w1505,w1504,w1503,w1502,w1501,w1500,w1499,w1498,w1497,w1496,w1495,w1494,w1493,w1492,w1491,w1490,w1489,w1488,w1487,w1486,w1485,w1484,w1483,w1482,w1481,w1480,w1479,w1478,w1477,w1476,w1475,w1474,w1473,w1472,w1471,w1470,w1469,w1468,w1467,w1466,w1465,w1464,w1463,w1462,w1461,w1460,w1459,w1458,w1457,w1456,w1455,w1454,w1453,w1452,w1451,w1450,w1449,w1448,w1447,w1446,w1445,w1444,w1443,w1442,w1441,w1440,w1439,w1438,w1437,w1436,w1435,w1434,w1433,w1432}, w1206, {w388,w387,w386,w385,w384,w383,w382,w381,w380,w379,w378,w377,w376,w375,w374,w373,w372,w371,w370,w369,w368,w367,w366,w365,w364,w363,w362,w361,w360,w359,w358,w357,w356,w355,w354,w353,w352,w351,w350,w349,w348,w347,w346,w345,w344,w343,w342,w341,w340,w339,w338,w337,w336,w335,w334,w333,w332,w331,w330,w329,w328,w327,w326,w325,w324,w323,w322,w321,w320,w319,w318,w317,w316,w315}, {w536,w535,w534,w533,w532,w531,w530,w529,w528,w527,w526,w525,w524,w523,w522,w521,w520,w519,w518,w517,w516,w515,w514,w513,w512,w511,w510,w509,w508,w507,w506,w505,w504,w503,w502,w501,w500,w499,w498,w497,w496,w495,w494,w493,w492,w491,w490,w489,w488,w487,w486,w485,w484,w483,w482,w481,w480,w479,w478,w477,w476,w475,w474,w473,w472,w471,w470,w469,w468,w467,w466,w465,w464,w463});
    wire w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284;
    sw_m #(.SIZE(74)) sw39({w3210,w3209,w3208,w3207,w3206,w3205,w3204,w3203,w3202,w3201,w3200,w3199,w3198,w3197,w3196,w3195,w3194,w3193,w3192,w3191,w3190,w3189,w3188,w3187,w3186,w3185,w3184,w3183,w3182,w3181,w3180,w3179,w3178,w3177,w3176,w3175,w3174,w3173,w3172,w3171,w3170,w3169,w3168,w3167,w3166,w3165,w3164,w3163,w3162,w3161,w3160,w3159,w3158,w3157,w3156,w3155,w3154,w3153,w3152,w3151,w3150,w3149,w3148,w3147,w3146,w3145,w3144,w3143,w3142,w3141,w3140,w3139,w3138,w3137}, {w3284,w3283,w3282,w3281,w3280,w3279,w3278,w3277,w3276,w3275,w3274,w3273,w3272,w3271,w3270,w3269,w3268,w3267,w3266,w3265,w3264,w3263,w3262,w3261,w3260,w3259,w3258,w3257,w3256,w3255,w3254,w3253,w3252,w3251,w3250,w3249,w3248,w3247,w3246,w3245,w3244,w3243,w3242,w3241,w3240,w3239,w3238,w3237,w3236,w3235,w3234,w3233,w3232,w3231,w3230,w3229,w3228,w3227,w3226,w3225,w3224,w3223,w3222,w3221,w3220,w3219,w3218,w3217,w3216,w3215,w3214,w3213,w3212,w3211}, w2985, {w462,w461,w460,w459,w458,w457,w456,w455,w454,w453,w452,w451,w450,w449,w448,w447,w446,w445,w444,w443,w442,w441,w440,w439,w438,w437,w436,w435,w434,w433,w432,w431,w430,w429,w428,w427,w426,w425,w424,w423,w422,w421,w420,w419,w418,w417,w416,w415,w414,w413,w412,w411,w410,w409,w408,w407,w406,w405,w404,w403,w402,w401,w400,w399,w398,w397,w396,w395,w394,w393,w392,w391,w390,w389}, {w610,w609,w608,w607,w606,w605,w604,w603,w602,w601,w600,w599,w598,w597,w596,w595,w594,w593,w592,w591,w590,w589,w588,w587,w586,w585,w584,w583,w582,w581,w580,w579,w578,w577,w576,w575,w574,w573,w572,w571,w570,w569,w568,w567,w566,w565,w564,w563,w562,w561,w560,w559,w558,w557,w556,w555,w554,w553,w552,w551,w550,w549,w548,w547,w546,w545,w544,w543,w542,w541,w540,w539,w538,w537});
    wire w1207;
    xor xor40(w1207, w1204, w1205);
    wire w2986;
    xor xor41(w2986, w2983, w2984);
    wire w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653;
    sw_m #(.SIZE(74)) sw42({w1579,w1578,w1577,w1576,w1575,w1574,w1573,w1572,w1571,w1570,w1569,w1568,w1567,w1566,w1565,w1564,w1563,w1562,w1561,w1560,w1559,w1558,w1557,w1556,w1555,w1554,w1553,w1552,w1551,w1550,w1549,w1548,w1547,w1546,w1545,w1544,w1543,w1542,w1541,w1540,w1539,w1538,w1537,w1536,w1535,w1534,w1533,w1532,w1531,w1530,w1529,w1528,w1527,w1526,w1525,w1524,w1523,w1522,w1521,w1520,w1519,w1518,w1517,w1516,w1515,w1514,w1513,w1512,w1511,w1510,w1509,w1508,w1507,w1506}, {w1653,w1652,w1651,w1650,w1649,w1648,w1647,w1646,w1645,w1644,w1643,w1642,w1641,w1640,w1639,w1638,w1637,w1636,w1635,w1634,w1633,w1632,w1631,w1630,w1629,w1628,w1627,w1626,w1625,w1624,w1623,w1622,w1621,w1620,w1619,w1618,w1617,w1616,w1615,w1614,w1613,w1612,w1611,w1610,w1609,w1608,w1607,w1606,w1605,w1604,w1603,w1602,w1601,w1600,w1599,w1598,w1597,w1596,w1595,w1594,w1593,w1592,w1591,w1590,w1589,w1588,w1587,w1586,w1585,w1584,w1583,w1582,w1581,w1580}, w1209, {w684,w683,w682,w681,w680,w679,w678,w677,w676,w675,w674,w673,w672,w671,w670,w669,w668,w667,w666,w665,w664,w663,w662,w661,w660,w659,w658,w657,w656,w655,w654,w653,w652,w651,w650,w649,w648,w647,w646,w645,w644,w643,w642,w641,w640,w639,w638,w637,w636,w635,w634,w633,w632,w631,w630,w629,w628,w627,w626,w625,w624,w623,w622,w621,w620,w619,w618,w617,w616,w615,w614,w613,w612,w611}, {w832,w831,w830,w829,w828,w827,w826,w825,w824,w823,w822,w821,w820,w819,w818,w817,w816,w815,w814,w813,w812,w811,w810,w809,w808,w807,w806,w805,w804,w803,w802,w801,w800,w799,w798,w797,w796,w795,w794,w793,w792,w791,w790,w789,w788,w787,w786,w785,w784,w783,w782,w781,w780,w779,w778,w777,w776,w775,w774,w773,w772,w771,w770,w769,w768,w767,w766,w765,w764,w763,w762,w761,w760,w759});
    wire w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951;
    sw_m #(.SIZE(74)) sw43({w1877,w1876,w1875,w1874,w1873,w1872,w1871,w1870,w1869,w1868,w1867,w1866,w1865,w1864,w1863,w1862,w1861,w1860,w1859,w1858,w1857,w1856,w1855,w1854,w1853,w1852,w1851,w1850,w1849,w1848,w1847,w1846,w1845,w1844,w1843,w1842,w1841,w1840,w1839,w1838,w1837,w1836,w1835,w1834,w1833,w1832,w1831,w1830,w1829,w1828,w1827,w1826,w1825,w1824,w1823,w1822,w1821,w1820,w1819,w1818,w1817,w1816,w1815,w1814,w1813,w1812,w1811,w1810,w1809,w1808,w1807,w1806,w1805,w1804}, {w1951,w1950,w1949,w1948,w1947,w1946,w1945,w1944,w1943,w1942,w1941,w1940,w1939,w1938,w1937,w1936,w1935,w1934,w1933,w1932,w1931,w1930,w1929,w1928,w1927,w1926,w1925,w1924,w1923,w1922,w1921,w1920,w1919,w1918,w1917,w1916,w1915,w1914,w1913,w1912,w1911,w1910,w1909,w1908,w1907,w1906,w1905,w1904,w1903,w1902,w1901,w1900,w1899,w1898,w1897,w1896,w1895,w1894,w1893,w1892,w1891,w1890,w1889,w1888,w1887,w1886,w1885,w1884,w1883,w1882,w1881,w1880,w1879,w1878}, w1283, {w1283,w1282,w1281,w1280,w1279,w1278,w1277,w1276,w1275,w1274,w1273,w1272,w1271,w1270,w1269,w1268,w1267,w1266,w1265,w1264,w1263,w1262,w1261,w1260,w1259,w1258,w1257,w1256,w1255,w1254,w1253,w1252,w1251,w1250,w1249,w1248,w1247,w1246,w1245,w1244,w1243,w1242,w1241,w1240,w1239,w1238,w1237,w1236,w1235,w1234,w1233,w1232,w1231,w1230,w1229,w1228,w1227,w1226,w1225,w1224,w1223,w1222,w1221,w1220,w1219,w1218,w1217,w1216,w1215,w1214,w1213,w1212,w1211,w1210}, {w1431,w1430,w1429,w1428,w1427,w1426,w1425,w1424,w1423,w1422,w1421,w1420,w1419,w1418,w1417,w1416,w1415,w1414,w1413,w1412,w1411,w1410,w1409,w1408,w1407,w1406,w1405,w1404,w1403,w1402,w1401,w1400,w1399,w1398,w1397,w1396,w1395,w1394,w1393,w1392,w1391,w1390,w1389,w1388,w1387,w1386,w1385,w1384,w1383,w1382,w1381,w1380,w1379,w1378,w1377,w1376,w1375,w1374,w1373,w1372,w1371,w1370,w1369,w1368,w1367,w1366,w1365,w1364,w1363,w1362,w1361,w1360,w1359,w1358});
    wire w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541;
    sw_m #(.SIZE(74)) sw44({w2467,w2466,w2465,w2464,w2463,w2462,w2461,w2460,w2459,w2458,w2457,w2456,w2455,w2454,w2453,w2452,w2451,w2450,w2449,w2448,w2447,w2446,w2445,w2444,w2443,w2442,w2441,w2440,w2439,w2438,w2437,w2436,w2435,w2434,w2433,w2432,w2431,w2430,w2429,w2428,w2427,w2426,w2425,w2424,w2423,w2422,w2421,w2420,w2419,w2418,w2417,w2416,w2415,w2414,w2413,w2412,w2411,w2410,w2409,w2408,w2407,w2406,w2405,w2404,w2403,w2402,w2401,w2400,w2399,w2398,w2397,w2396,w2395,w2394}, {w2541,w2540,w2539,w2538,w2537,w2536,w2535,w2534,w2533,w2532,w2531,w2530,w2529,w2528,w2527,w2526,w2525,w2524,w2523,w2522,w2521,w2520,w2519,w2518,w2517,w2516,w2515,w2514,w2513,w2512,w2511,w2510,w2509,w2508,w2507,w2506,w2505,w2504,w2503,w2502,w2501,w2500,w2499,w2498,w2497,w2496,w2495,w2494,w2493,w2492,w2491,w2490,w2489,w2488,w2487,w2486,w2485,w2484,w2483,w2482,w2481,w2480,w2479,w2478,w2477,w2476,w2475,w2474,w2473,w2472,w2471,w2470,w2469,w2468}, w1357, {w1357,w1356,w1355,w1354,w1353,w1352,w1351,w1350,w1349,w1348,w1347,w1346,w1345,w1344,w1343,w1342,w1341,w1340,w1339,w1338,w1337,w1336,w1335,w1334,w1333,w1332,w1331,w1330,w1329,w1328,w1327,w1326,w1325,w1324,w1323,w1322,w1321,w1320,w1319,w1318,w1317,w1316,w1315,w1314,w1313,w1312,w1311,w1310,w1309,w1308,w1307,w1306,w1305,w1304,w1303,w1302,w1301,w1300,w1299,w1298,w1297,w1296,w1295,w1294,w1293,w1292,w1291,w1290,w1289,w1288,w1287,w1286,w1285,w1284}, {w1505,w1504,w1503,w1502,w1501,w1500,w1499,w1498,w1497,w1496,w1495,w1494,w1493,w1492,w1491,w1490,w1489,w1488,w1487,w1486,w1485,w1484,w1483,w1482,w1481,w1480,w1479,w1478,w1477,w1476,w1475,w1474,w1473,w1472,w1471,w1470,w1469,w1468,w1467,w1466,w1465,w1464,w1463,w1462,w1461,w1460,w1459,w1458,w1457,w1456,w1455,w1454,w1453,w1452,w1451,w1450,w1449,w1448,w1447,w1446,w1445,w1444,w1443,w1442,w1441,w1440,w1439,w1438,w1437,w1436,w1435,w1434,w1433,w1432});
    wire w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432;
    sw_m #(.SIZE(74)) sw45({w3358,w3357,w3356,w3355,w3354,w3353,w3352,w3351,w3350,w3349,w3348,w3347,w3346,w3345,w3344,w3343,w3342,w3341,w3340,w3339,w3338,w3337,w3336,w3335,w3334,w3333,w3332,w3331,w3330,w3329,w3328,w3327,w3326,w3325,w3324,w3323,w3322,w3321,w3320,w3319,w3318,w3317,w3316,w3315,w3314,w3313,w3312,w3311,w3310,w3309,w3308,w3307,w3306,w3305,w3304,w3303,w3302,w3301,w3300,w3299,w3298,w3297,w3296,w3295,w3294,w3293,w3292,w3291,w3290,w3289,w3288,w3287,w3286,w3285}, {w3432,w3431,w3430,w3429,w3428,w3427,w3426,w3425,w3424,w3423,w3422,w3421,w3420,w3419,w3418,w3417,w3416,w3415,w3414,w3413,w3412,w3411,w3410,w3409,w3408,w3407,w3406,w3405,w3404,w3403,w3402,w3401,w3400,w3399,w3398,w3397,w3396,w3395,w3394,w3393,w3392,w3391,w3390,w3389,w3388,w3387,w3386,w3385,w3384,w3383,w3382,w3381,w3380,w3379,w3378,w3377,w3376,w3375,w3374,w3373,w3372,w3371,w3370,w3369,w3368,w3367,w3366,w3365,w3364,w3363,w3362,w3361,w3360,w3359}, w2988, {w758,w757,w756,w755,w754,w753,w752,w751,w750,w749,w748,w747,w746,w745,w744,w743,w742,w741,w740,w739,w738,w737,w736,w735,w734,w733,w732,w731,w730,w729,w728,w727,w726,w725,w724,w723,w722,w721,w720,w719,w718,w717,w716,w715,w714,w713,w712,w711,w710,w709,w708,w707,w706,w705,w704,w703,w702,w701,w700,w699,w698,w697,w696,w695,w694,w693,w692,w691,w690,w689,w688,w687,w686,w685}, {w906,w905,w904,w903,w902,w901,w900,w899,w898,w897,w896,w895,w894,w893,w892,w891,w890,w889,w888,w887,w886,w885,w884,w883,w882,w881,w880,w879,w878,w877,w876,w875,w874,w873,w872,w871,w870,w869,w868,w867,w866,w865,w864,w863,w862,w861,w860,w859,w858,w857,w856,w855,w854,w853,w852,w851,w850,w849,w848,w847,w846,w845,w844,w843,w842,w841,w840,w839,w838,w837,w836,w835,w834,w833});
    wire w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730;
    sw_m #(.SIZE(74)) sw46({w3656,w3655,w3654,w3653,w3652,w3651,w3650,w3649,w3648,w3647,w3646,w3645,w3644,w3643,w3642,w3641,w3640,w3639,w3638,w3637,w3636,w3635,w3634,w3633,w3632,w3631,w3630,w3629,w3628,w3627,w3626,w3625,w3624,w3623,w3622,w3621,w3620,w3619,w3618,w3617,w3616,w3615,w3614,w3613,w3612,w3611,w3610,w3609,w3608,w3607,w3606,w3605,w3604,w3603,w3602,w3601,w3600,w3599,w3598,w3597,w3596,w3595,w3594,w3593,w3592,w3591,w3590,w3589,w3588,w3587,w3586,w3585,w3584,w3583}, {w3730,w3729,w3728,w3727,w3726,w3725,w3724,w3723,w3722,w3721,w3720,w3719,w3718,w3717,w3716,w3715,w3714,w3713,w3712,w3711,w3710,w3709,w3708,w3707,w3706,w3705,w3704,w3703,w3702,w3701,w3700,w3699,w3698,w3697,w3696,w3695,w3694,w3693,w3692,w3691,w3690,w3689,w3688,w3687,w3686,w3685,w3684,w3683,w3682,w3681,w3680,w3679,w3678,w3677,w3676,w3675,w3674,w3673,w3672,w3671,w3670,w3669,w3668,w3667,w3666,w3665,w3664,w3663,w3662,w3661,w3660,w3659,w3658,w3657}, w3062, {w3062,w3061,w3060,w3059,w3058,w3057,w3056,w3055,w3054,w3053,w3052,w3051,w3050,w3049,w3048,w3047,w3046,w3045,w3044,w3043,w3042,w3041,w3040,w3039,w3038,w3037,w3036,w3035,w3034,w3033,w3032,w3031,w3030,w3029,w3028,w3027,w3026,w3025,w3024,w3023,w3022,w3021,w3020,w3019,w3018,w3017,w3016,w3015,w3014,w3013,w3012,w3011,w3010,w3009,w3008,w3007,w3006,w3005,w3004,w3003,w3002,w3001,w3000,w2999,w2998,w2997,w2996,w2995,w2994,w2993,w2992,w2991,w2990,w2989}, {w3210,w3209,w3208,w3207,w3206,w3205,w3204,w3203,w3202,w3201,w3200,w3199,w3198,w3197,w3196,w3195,w3194,w3193,w3192,w3191,w3190,w3189,w3188,w3187,w3186,w3185,w3184,w3183,w3182,w3181,w3180,w3179,w3178,w3177,w3176,w3175,w3174,w3173,w3172,w3171,w3170,w3169,w3168,w3167,w3166,w3165,w3164,w3163,w3162,w3161,w3160,w3159,w3158,w3157,w3156,w3155,w3154,w3153,w3152,w3151,w3150,w3149,w3148,w3147,w3146,w3145,w3144,w3143,w3142,w3141,w3140,w3139,w3138,w3137});
    wire w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320;
    sw_m #(.SIZE(74)) sw47({w4246,w4245,w4244,w4243,w4242,w4241,w4240,w4239,w4238,w4237,w4236,w4235,w4234,w4233,w4232,w4231,w4230,w4229,w4228,w4227,w4226,w4225,w4224,w4223,w4222,w4221,w4220,w4219,w4218,w4217,w4216,w4215,w4214,w4213,w4212,w4211,w4210,w4209,w4208,w4207,w4206,w4205,w4204,w4203,w4202,w4201,w4200,w4199,w4198,w4197,w4196,w4195,w4194,w4193,w4192,w4191,w4190,w4189,w4188,w4187,w4186,w4185,w4184,w4183,w4182,w4181,w4180,w4179,w4178,w4177,w4176,w4175,w4174,w4173}, {w4320,w4319,w4318,w4317,w4316,w4315,w4314,w4313,w4312,w4311,w4310,w4309,w4308,w4307,w4306,w4305,w4304,w4303,w4302,w4301,w4300,w4299,w4298,w4297,w4296,w4295,w4294,w4293,w4292,w4291,w4290,w4289,w4288,w4287,w4286,w4285,w4284,w4283,w4282,w4281,w4280,w4279,w4278,w4277,w4276,w4275,w4274,w4273,w4272,w4271,w4270,w4269,w4268,w4267,w4266,w4265,w4264,w4263,w4262,w4261,w4260,w4259,w4258,w4257,w4256,w4255,w4254,w4253,w4252,w4251,w4250,w4249,w4248,w4247}, w3136, {w3136,w3135,w3134,w3133,w3132,w3131,w3130,w3129,w3128,w3127,w3126,w3125,w3124,w3123,w3122,w3121,w3120,w3119,w3118,w3117,w3116,w3115,w3114,w3113,w3112,w3111,w3110,w3109,w3108,w3107,w3106,w3105,w3104,w3103,w3102,w3101,w3100,w3099,w3098,w3097,w3096,w3095,w3094,w3093,w3092,w3091,w3090,w3089,w3088,w3087,w3086,w3085,w3084,w3083,w3082,w3081,w3080,w3079,w3078,w3077,w3076,w3075,w3074,w3073,w3072,w3071,w3070,w3069,w3068,w3067,w3066,w3065,w3064,w3063}, {w3284,w3283,w3282,w3281,w3280,w3279,w3278,w3277,w3276,w3275,w3274,w3273,w3272,w3271,w3270,w3269,w3268,w3267,w3266,w3265,w3264,w3263,w3262,w3261,w3260,w3259,w3258,w3257,w3256,w3255,w3254,w3253,w3252,w3251,w3250,w3249,w3248,w3247,w3246,w3245,w3244,w3243,w3242,w3241,w3240,w3239,w3238,w3237,w3236,w3235,w3234,w3233,w3232,w3231,w3230,w3229,w3228,w3227,w3226,w3225,w3224,w3223,w3222,w3221,w3220,w3219,w3218,w3217,w3216,w3215,w3214,w3213,w3212,w3211});
    wire w1208;
    xor xor48(w1208, w1206, w1207);
    wire w1802;
    xor xor49(w1802, w1431, w1579);
    wire w2392;
    xor xor50(w2392, w1505, w1653);
    wire w2987;
    xor xor51(w2987, w2985, w2986);
    wire w3581;
    xor xor52(w3581, w3210, w3358);
    wire w4171;
    xor xor53(w4171, w3284, w3432);
    wire w1803;
    xor xor54(w1803, w1283, w1802);
    wire w2393;
    xor xor55(w2393, w1357, w2392);
    wire w3582;
    xor xor56(w3582, w3062, w3581);
    wire w4172;
    xor xor57(w4172, w3136, w4171);
    wire w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801;
    sw_m #(.SIZE(74)) sw58({w1727,w1726,w1725,w1724,w1723,w1722,w1721,w1720,w1719,w1718,w1717,w1716,w1715,w1714,w1713,w1712,w1711,w1710,w1709,w1708,w1707,w1706,w1705,w1704,w1703,w1702,w1701,w1700,w1699,w1698,w1697,w1696,w1695,w1694,w1693,w1692,w1691,w1690,w1689,w1688,w1687,w1686,w1685,w1684,w1683,w1682,w1681,w1680,w1679,w1678,w1677,w1676,w1675,w1674,w1673,w1672,w1671,w1670,w1669,w1668,w1667,w1666,w1665,w1664,w1663,w1662,w1661,w1660,w1659,w1658,w1657,w1656,w1655,w1654}, {w1801,w1800,w1799,w1798,w1797,w1796,w1795,w1794,w1793,w1792,w1791,w1790,w1789,w1788,w1787,w1786,w1785,w1784,w1783,w1782,w1781,w1780,w1779,w1778,w1777,w1776,w1775,w1774,w1773,w1772,w1771,w1770,w1769,w1768,w1767,w1766,w1765,w1764,w1763,w1762,w1761,w1760,w1759,w1758,w1757,w1756,w1755,w1754,w1753,w1752,w1751,w1750,w1749,w1748,w1747,w1746,w1745,w1744,w1743,w1742,w1741,w1740,w1739,w1738,w1737,w1736,w1735,w1734,w1733,w1732,w1731,w1730,w1729,w1728}, w1208, {w980,w979,w978,w977,w976,w975,w974,w973,w972,w971,w970,w969,w968,w967,w966,w965,w964,w963,w962,w961,w960,w959,w958,w957,w956,w955,w954,w953,w952,w951,w950,w949,w948,w947,w946,w945,w944,w943,w942,w941,w940,w939,w938,w937,w936,w935,w934,w933,w932,w931,w930,w929,w928,w927,w926,w925,w924,w923,w922,w921,w920,w919,w918,w917,w916,w915,w914,w913,w912,w911,w910,w909,w908,w907}, {w1128,w1127,w1126,w1125,w1124,w1123,w1122,w1121,w1120,w1119,w1118,w1117,w1116,w1115,w1114,w1113,w1112,w1111,w1110,w1109,w1108,w1107,w1106,w1105,w1104,w1103,w1102,w1101,w1100,w1099,w1098,w1097,w1096,w1095,w1094,w1093,w1092,w1091,w1090,w1089,w1088,w1087,w1086,w1085,w1084,w1083,w1082,w1081,w1080,w1079,w1078,w1077,w1076,w1075,w1074,w1073,w1072,w1071,w1070,w1069,w1068,w1067,w1066,w1065,w1064,w1063,w1062,w1061,w1060,w1059,w1058,w1057,w1056,w1055});
    wire w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580;
    sw_m #(.SIZE(74)) sw59({w3506,w3505,w3504,w3503,w3502,w3501,w3500,w3499,w3498,w3497,w3496,w3495,w3494,w3493,w3492,w3491,w3490,w3489,w3488,w3487,w3486,w3485,w3484,w3483,w3482,w3481,w3480,w3479,w3478,w3477,w3476,w3475,w3474,w3473,w3472,w3471,w3470,w3469,w3468,w3467,w3466,w3465,w3464,w3463,w3462,w3461,w3460,w3459,w3458,w3457,w3456,w3455,w3454,w3453,w3452,w3451,w3450,w3449,w3448,w3447,w3446,w3445,w3444,w3443,w3442,w3441,w3440,w3439,w3438,w3437,w3436,w3435,w3434,w3433}, {w3580,w3579,w3578,w3577,w3576,w3575,w3574,w3573,w3572,w3571,w3570,w3569,w3568,w3567,w3566,w3565,w3564,w3563,w3562,w3561,w3560,w3559,w3558,w3557,w3556,w3555,w3554,w3553,w3552,w3551,w3550,w3549,w3548,w3547,w3546,w3545,w3544,w3543,w3542,w3541,w3540,w3539,w3538,w3537,w3536,w3535,w3534,w3533,w3532,w3531,w3530,w3529,w3528,w3527,w3526,w3525,w3524,w3523,w3522,w3521,w3520,w3519,w3518,w3517,w3516,w3515,w3514,w3513,w3512,w3511,w3510,w3509,w3508,w3507}, w2987, {w1054,w1053,w1052,w1051,w1050,w1049,w1048,w1047,w1046,w1045,w1044,w1043,w1042,w1041,w1040,w1039,w1038,w1037,w1036,w1035,w1034,w1033,w1032,w1031,w1030,w1029,w1028,w1027,w1026,w1025,w1024,w1023,w1022,w1021,w1020,w1019,w1018,w1017,w1016,w1015,w1014,w1013,w1012,w1011,w1010,w1009,w1008,w1007,w1006,w1005,w1004,w1003,w1002,w1001,w1000,w999,w998,w997,w996,w995,w994,w993,w992,w991,w990,w989,w988,w987,w986,w985,w984,w983,w982,w981}, {w1202,w1201,w1200,w1199,w1198,w1197,w1196,w1195,w1194,w1193,w1192,w1191,w1190,w1189,w1188,w1187,w1186,w1185,w1184,w1183,w1182,w1181,w1180,w1179,w1178,w1177,w1176,w1175,w1174,w1173,w1172,w1171,w1170,w1169,w1168,w1167,w1166,w1165,w1164,w1163,w1162,w1161,w1160,w1159,w1158,w1157,w1156,w1155,w1154,w1153,w1152,w1151,w1150,w1149,w1148,w1147,w1146,w1145,w1144,w1143,w1142,w1141,w1140,w1139,w1138,w1137,w1136,w1135,w1134,w1133,w1132,w1131,w1130,w1129});
    wire w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099;
    sw_m #(.SIZE(74)) sw60({w2025,w2024,w2023,w2022,w2021,w2020,w2019,w2018,w2017,w2016,w2015,w2014,w2013,w2012,w2011,w2010,w2009,w2008,w2007,w2006,w2005,w2004,w2003,w2002,w2001,w2000,w1999,w1998,w1997,w1996,w1995,w1994,w1993,w1992,w1991,w1990,w1989,w1988,w1987,w1986,w1985,w1984,w1983,w1982,w1981,w1980,w1979,w1978,w1977,w1976,w1975,w1974,w1973,w1972,w1971,w1970,w1969,w1968,w1967,w1966,w1965,w1964,w1963,w1962,w1961,w1960,w1959,w1958,w1957,w1956,w1955,w1954,w1953,w1952}, {w2099,w2098,w2097,w2096,w2095,w2094,w2093,w2092,w2091,w2090,w2089,w2088,w2087,w2086,w2085,w2084,w2083,w2082,w2081,w2080,w2079,w2078,w2077,w2076,w2075,w2074,w2073,w2072,w2071,w2070,w2069,w2068,w2067,w2066,w2065,w2064,w2063,w2062,w2061,w2060,w2059,w2058,w2057,w2056,w2055,w2054,w2053,w2052,w2051,w2050,w2049,w2048,w2047,w2046,w2045,w2044,w2043,w2042,w2041,w2040,w2039,w2038,w2037,w2036,w2035,w2034,w2033,w2032,w2031,w2030,w2029,w2028,w2027,w2026}, w1803, {w1579,w1578,w1577,w1576,w1575,w1574,w1573,w1572,w1571,w1570,w1569,w1568,w1567,w1566,w1565,w1564,w1563,w1562,w1561,w1560,w1559,w1558,w1557,w1556,w1555,w1554,w1553,w1552,w1551,w1550,w1549,w1548,w1547,w1546,w1545,w1544,w1543,w1542,w1541,w1540,w1539,w1538,w1537,w1536,w1535,w1534,w1533,w1532,w1531,w1530,w1529,w1528,w1527,w1526,w1525,w1524,w1523,w1522,w1521,w1520,w1519,w1518,w1517,w1516,w1515,w1514,w1513,w1512,w1511,w1510,w1509,w1508,w1507,w1506}, {w1727,w1726,w1725,w1724,w1723,w1722,w1721,w1720,w1719,w1718,w1717,w1716,w1715,w1714,w1713,w1712,w1711,w1710,w1709,w1708,w1707,w1706,w1705,w1704,w1703,w1702,w1701,w1700,w1699,w1698,w1697,w1696,w1695,w1694,w1693,w1692,w1691,w1690,w1689,w1688,w1687,w1686,w1685,w1684,w1683,w1682,w1681,w1680,w1679,w1678,w1677,w1676,w1675,w1674,w1673,w1672,w1671,w1670,w1669,w1668,w1667,w1666,w1665,w1664,w1663,w1662,w1661,w1660,w1659,w1658,w1657,w1656,w1655,w1654});
    wire w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689;
    sw_m #(.SIZE(74)) sw61({w2615,w2614,w2613,w2612,w2611,w2610,w2609,w2608,w2607,w2606,w2605,w2604,w2603,w2602,w2601,w2600,w2599,w2598,w2597,w2596,w2595,w2594,w2593,w2592,w2591,w2590,w2589,w2588,w2587,w2586,w2585,w2584,w2583,w2582,w2581,w2580,w2579,w2578,w2577,w2576,w2575,w2574,w2573,w2572,w2571,w2570,w2569,w2568,w2567,w2566,w2565,w2564,w2563,w2562,w2561,w2560,w2559,w2558,w2557,w2556,w2555,w2554,w2553,w2552,w2551,w2550,w2549,w2548,w2547,w2546,w2545,w2544,w2543,w2542}, {w2689,w2688,w2687,w2686,w2685,w2684,w2683,w2682,w2681,w2680,w2679,w2678,w2677,w2676,w2675,w2674,w2673,w2672,w2671,w2670,w2669,w2668,w2667,w2666,w2665,w2664,w2663,w2662,w2661,w2660,w2659,w2658,w2657,w2656,w2655,w2654,w2653,w2652,w2651,w2650,w2649,w2648,w2647,w2646,w2645,w2644,w2643,w2642,w2641,w2640,w2639,w2638,w2637,w2636,w2635,w2634,w2633,w2632,w2631,w2630,w2629,w2628,w2627,w2626,w2625,w2624,w2623,w2622,w2621,w2620,w2619,w2618,w2617,w2616}, w2393, {w1653,w1652,w1651,w1650,w1649,w1648,w1647,w1646,w1645,w1644,w1643,w1642,w1641,w1640,w1639,w1638,w1637,w1636,w1635,w1634,w1633,w1632,w1631,w1630,w1629,w1628,w1627,w1626,w1625,w1624,w1623,w1622,w1621,w1620,w1619,w1618,w1617,w1616,w1615,w1614,w1613,w1612,w1611,w1610,w1609,w1608,w1607,w1606,w1605,w1604,w1603,w1602,w1601,w1600,w1599,w1598,w1597,w1596,w1595,w1594,w1593,w1592,w1591,w1590,w1589,w1588,w1587,w1586,w1585,w1584,w1583,w1582,w1581,w1580}, {w1801,w1800,w1799,w1798,w1797,w1796,w1795,w1794,w1793,w1792,w1791,w1790,w1789,w1788,w1787,w1786,w1785,w1784,w1783,w1782,w1781,w1780,w1779,w1778,w1777,w1776,w1775,w1774,w1773,w1772,w1771,w1770,w1769,w1768,w1767,w1766,w1765,w1764,w1763,w1762,w1761,w1760,w1759,w1758,w1757,w1756,w1755,w1754,w1753,w1752,w1751,w1750,w1749,w1748,w1747,w1746,w1745,w1744,w1743,w1742,w1741,w1740,w1739,w1738,w1737,w1736,w1735,w1734,w1733,w1732,w1731,w1730,w1729,w1728});
    wire w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878;
    sw_m #(.SIZE(74)) sw62({w3804,w3803,w3802,w3801,w3800,w3799,w3798,w3797,w3796,w3795,w3794,w3793,w3792,w3791,w3790,w3789,w3788,w3787,w3786,w3785,w3784,w3783,w3782,w3781,w3780,w3779,w3778,w3777,w3776,w3775,w3774,w3773,w3772,w3771,w3770,w3769,w3768,w3767,w3766,w3765,w3764,w3763,w3762,w3761,w3760,w3759,w3758,w3757,w3756,w3755,w3754,w3753,w3752,w3751,w3750,w3749,w3748,w3747,w3746,w3745,w3744,w3743,w3742,w3741,w3740,w3739,w3738,w3737,w3736,w3735,w3734,w3733,w3732,w3731}, {w3878,w3877,w3876,w3875,w3874,w3873,w3872,w3871,w3870,w3869,w3868,w3867,w3866,w3865,w3864,w3863,w3862,w3861,w3860,w3859,w3858,w3857,w3856,w3855,w3854,w3853,w3852,w3851,w3850,w3849,w3848,w3847,w3846,w3845,w3844,w3843,w3842,w3841,w3840,w3839,w3838,w3837,w3836,w3835,w3834,w3833,w3832,w3831,w3830,w3829,w3828,w3827,w3826,w3825,w3824,w3823,w3822,w3821,w3820,w3819,w3818,w3817,w3816,w3815,w3814,w3813,w3812,w3811,w3810,w3809,w3808,w3807,w3806,w3805}, w3582, {w3358,w3357,w3356,w3355,w3354,w3353,w3352,w3351,w3350,w3349,w3348,w3347,w3346,w3345,w3344,w3343,w3342,w3341,w3340,w3339,w3338,w3337,w3336,w3335,w3334,w3333,w3332,w3331,w3330,w3329,w3328,w3327,w3326,w3325,w3324,w3323,w3322,w3321,w3320,w3319,w3318,w3317,w3316,w3315,w3314,w3313,w3312,w3311,w3310,w3309,w3308,w3307,w3306,w3305,w3304,w3303,w3302,w3301,w3300,w3299,w3298,w3297,w3296,w3295,w3294,w3293,w3292,w3291,w3290,w3289,w3288,w3287,w3286,w3285}, {w3506,w3505,w3504,w3503,w3502,w3501,w3500,w3499,w3498,w3497,w3496,w3495,w3494,w3493,w3492,w3491,w3490,w3489,w3488,w3487,w3486,w3485,w3484,w3483,w3482,w3481,w3480,w3479,w3478,w3477,w3476,w3475,w3474,w3473,w3472,w3471,w3470,w3469,w3468,w3467,w3466,w3465,w3464,w3463,w3462,w3461,w3460,w3459,w3458,w3457,w3456,w3455,w3454,w3453,w3452,w3451,w3450,w3449,w3448,w3447,w3446,w3445,w3444,w3443,w3442,w3441,w3440,w3439,w3438,w3437,w3436,w3435,w3434,w3433});
    wire w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468;
    sw_m #(.SIZE(74)) sw63({w4394,w4393,w4392,w4391,w4390,w4389,w4388,w4387,w4386,w4385,w4384,w4383,w4382,w4381,w4380,w4379,w4378,w4377,w4376,w4375,w4374,w4373,w4372,w4371,w4370,w4369,w4368,w4367,w4366,w4365,w4364,w4363,w4362,w4361,w4360,w4359,w4358,w4357,w4356,w4355,w4354,w4353,w4352,w4351,w4350,w4349,w4348,w4347,w4346,w4345,w4344,w4343,w4342,w4341,w4340,w4339,w4338,w4337,w4336,w4335,w4334,w4333,w4332,w4331,w4330,w4329,w4328,w4327,w4326,w4325,w4324,w4323,w4322,w4321}, {w4468,w4467,w4466,w4465,w4464,w4463,w4462,w4461,w4460,w4459,w4458,w4457,w4456,w4455,w4454,w4453,w4452,w4451,w4450,w4449,w4448,w4447,w4446,w4445,w4444,w4443,w4442,w4441,w4440,w4439,w4438,w4437,w4436,w4435,w4434,w4433,w4432,w4431,w4430,w4429,w4428,w4427,w4426,w4425,w4424,w4423,w4422,w4421,w4420,w4419,w4418,w4417,w4416,w4415,w4414,w4413,w4412,w4411,w4410,w4409,w4408,w4407,w4406,w4405,w4404,w4403,w4402,w4401,w4400,w4399,w4398,w4397,w4396,w4395}, w4172, {w3432,w3431,w3430,w3429,w3428,w3427,w3426,w3425,w3424,w3423,w3422,w3421,w3420,w3419,w3418,w3417,w3416,w3415,w3414,w3413,w3412,w3411,w3410,w3409,w3408,w3407,w3406,w3405,w3404,w3403,w3402,w3401,w3400,w3399,w3398,w3397,w3396,w3395,w3394,w3393,w3392,w3391,w3390,w3389,w3388,w3387,w3386,w3385,w3384,w3383,w3382,w3381,w3380,w3379,w3378,w3377,w3376,w3375,w3374,w3373,w3372,w3371,w3370,w3369,w3368,w3367,w3366,w3365,w3364,w3363,w3362,w3361,w3360,w3359}, {w3580,w3579,w3578,w3577,w3576,w3575,w3574,w3573,w3572,w3571,w3570,w3569,w3568,w3567,w3566,w3565,w3564,w3563,w3562,w3561,w3560,w3559,w3558,w3557,w3556,w3555,w3554,w3553,w3552,w3551,w3550,w3549,w3548,w3547,w3546,w3545,w3544,w3543,w3542,w3541,w3540,w3539,w3538,w3537,w3536,w3535,w3534,w3533,w3532,w3531,w3530,w3529,w3528,w3527,w3526,w3525,w3524,w3523,w3522,w3521,w3520,w3519,w3518,w3517,w3516,w3515,w3514,w3513,w3512,w3511,w3510,w3509,w3508,w3507});
    wire w2169, w2170, w2171, w2172, w2242, w2243, w2244, w2245;
    sw_m #(.SIZE(73)) sw64({w2172,w2171,w2170,w2169,w2168,w2167,w2166,w2165,w2164,w2163,w2162,w2161,w2160,w2159,w2158,w2157,w2156,w2155,w2154,w2153,w2152,w2151,w2150,w2149,w2148,w2147,w2146,w2145,w2144,w2143,w2142,w2141,w2140,w2139,w2138,w2137,w2136,w2135,w2134,w2133,w2132,w2131,w2130,w2129,w2128,w2127,w2126,w2125,w2124,w2123,w2122,w2121,w2120,w2119,w2118,w2117,w2116,w2115,w2114,w2113,w2112,w2111,w2110,w2109,w2108,w2107,w2106,w2105,w2104,w2103,w2102,w2101,w2100}, {w2245,w2244,w2243,w2242,w2241,w2240,w2239,w2238,w2237,w2236,w2235,w2234,w2233,w2232,w2231,w2230,w2229,w2228,w2227,w2226,w2225,w2224,w2223,w2222,w2221,w2220,w2219,w2218,w2217,w2216,w2215,w2214,w2213,w2212,w2211,w2210,w2209,w2208,w2207,w2206,w2205,w2204,w2203,w2202,w2201,w2200,w2199,w2198,w2197,w2196,w2195,w2194,w2193,w2192,w2191,w2190,w2189,w2188,w2187,w2186,w2185,w2184,w2183,w2182,w2181,w2180,w2179,w2178,w2177,w2176,w2175,w2174,w2173}, w1877, {w1876,w1875,w1874,w1873,w1872,w1871,w1870,w1869,w1868,w1867,w1866,w1865,w1864,w1863,w1862,w1861,w1860,w1859,w1858,w1857,w1856,w1855,w1854,w1853,w1852,w1851,w1850,w1849,w1848,w1847,w1846,w1845,w1844,w1843,w1842,w1841,w1840,w1839,w1838,w1837,w1836,w1835,w1834,w1833,w1832,w1831,w1830,w1829,w1828,w1827,w1826,w1825,w1824,w1823,w1822,w1821,w1820,w1819,w1818,w1817,w1816,w1815,w1814,w1813,w1812,w1811,w1810,w1809,w1808,w1807,w1806,w1805,w1804}, {w2024,w2023,w2022,w2021,w2020,w2019,w2018,w2017,w2016,w2015,w2014,w2013,w2012,w2011,w2010,w2009,w2008,w2007,w2006,w2005,w2004,w2003,w2002,w2001,w2000,w1999,w1998,w1997,w1996,w1995,w1994,w1993,w1992,w1991,w1990,w1989,w1988,w1987,w1986,w1985,w1984,w1983,w1982,w1981,w1980,w1979,w1978,w1977,w1976,w1975,w1974,w1973,w1972,w1971,w1970,w1969,w1968,w1967,w1966,w1965,w1964,w1963,w1962,w1961,w1960,w1959,w1958,w1957,w1956,w1955,w1954,w1953,w1952});
    wire w2315, w2316, w2317, w2318, w2388, w2389, w2390, w2391;
    sw_m #(.SIZE(73)) sw65({w2318,w2317,w2316,w2315,w2314,w2313,w2312,w2311,w2310,w2309,w2308,w2307,w2306,w2305,w2304,w2303,w2302,w2301,w2300,w2299,w2298,w2297,w2296,w2295,w2294,w2293,w2292,w2291,w2290,w2289,w2288,w2287,w2286,w2285,w2284,w2283,w2282,w2281,w2280,w2279,w2278,w2277,w2276,w2275,w2274,w2273,w2272,w2271,w2270,w2269,w2268,w2267,w2266,w2265,w2264,w2263,w2262,w2261,w2260,w2259,w2258,w2257,w2256,w2255,w2254,w2253,w2252,w2251,w2250,w2249,w2248,w2247,w2246}, {w2391,w2390,w2389,w2388,w2387,w2386,w2385,w2384,w2383,w2382,w2381,w2380,w2379,w2378,w2377,w2376,w2375,w2374,w2373,w2372,w2371,w2370,w2369,w2368,w2367,w2366,w2365,w2364,w2363,w2362,w2361,w2360,w2359,w2358,w2357,w2356,w2355,w2354,w2353,w2352,w2351,w2350,w2349,w2348,w2347,w2346,w2345,w2344,w2343,w2342,w2341,w2340,w2339,w2338,w2337,w2336,w2335,w2334,w2333,w2332,w2331,w2330,w2329,w2328,w2327,w2326,w2325,w2324,w2323,w2322,w2321,w2320,w2319}, w1951, {w1950,w1949,w1948,w1947,w1946,w1945,w1944,w1943,w1942,w1941,w1940,w1939,w1938,w1937,w1936,w1935,w1934,w1933,w1932,w1931,w1930,w1929,w1928,w1927,w1926,w1925,w1924,w1923,w1922,w1921,w1920,w1919,w1918,w1917,w1916,w1915,w1914,w1913,w1912,w1911,w1910,w1909,w1908,w1907,w1906,w1905,w1904,w1903,w1902,w1901,w1900,w1899,w1898,w1897,w1896,w1895,w1894,w1893,w1892,w1891,w1890,w1889,w1888,w1887,w1886,w1885,w1884,w1883,w1882,w1881,w1880,w1879,w1878}, {w2098,w2097,w2096,w2095,w2094,w2093,w2092,w2091,w2090,w2089,w2088,w2087,w2086,w2085,w2084,w2083,w2082,w2081,w2080,w2079,w2078,w2077,w2076,w2075,w2074,w2073,w2072,w2071,w2070,w2069,w2068,w2067,w2066,w2065,w2064,w2063,w2062,w2061,w2060,w2059,w2058,w2057,w2056,w2055,w2054,w2053,w2052,w2051,w2050,w2049,w2048,w2047,w2046,w2045,w2044,w2043,w2042,w2041,w2040,w2039,w2038,w2037,w2036,w2035,w2034,w2033,w2032,w2031,w2030,w2029,w2028,w2027,w2026});
    wire w2759, w2760, w2761, w2762, w2832, w2833, w2834, w2835;
    sw_m #(.SIZE(73)) sw66({w2762,w2761,w2760,w2759,w2758,w2757,w2756,w2755,w2754,w2753,w2752,w2751,w2750,w2749,w2748,w2747,w2746,w2745,w2744,w2743,w2742,w2741,w2740,w2739,w2738,w2737,w2736,w2735,w2734,w2733,w2732,w2731,w2730,w2729,w2728,w2727,w2726,w2725,w2724,w2723,w2722,w2721,w2720,w2719,w2718,w2717,w2716,w2715,w2714,w2713,w2712,w2711,w2710,w2709,w2708,w2707,w2706,w2705,w2704,w2703,w2702,w2701,w2700,w2699,w2698,w2697,w2696,w2695,w2694,w2693,w2692,w2691,w2690}, {w2835,w2834,w2833,w2832,w2831,w2830,w2829,w2828,w2827,w2826,w2825,w2824,w2823,w2822,w2821,w2820,w2819,w2818,w2817,w2816,w2815,w2814,w2813,w2812,w2811,w2810,w2809,w2808,w2807,w2806,w2805,w2804,w2803,w2802,w2801,w2800,w2799,w2798,w2797,w2796,w2795,w2794,w2793,w2792,w2791,w2790,w2789,w2788,w2787,w2786,w2785,w2784,w2783,w2782,w2781,w2780,w2779,w2778,w2777,w2776,w2775,w2774,w2773,w2772,w2771,w2770,w2769,w2768,w2767,w2766,w2765,w2764,w2763}, w2467, {w2466,w2465,w2464,w2463,w2462,w2461,w2460,w2459,w2458,w2457,w2456,w2455,w2454,w2453,w2452,w2451,w2450,w2449,w2448,w2447,w2446,w2445,w2444,w2443,w2442,w2441,w2440,w2439,w2438,w2437,w2436,w2435,w2434,w2433,w2432,w2431,w2430,w2429,w2428,w2427,w2426,w2425,w2424,w2423,w2422,w2421,w2420,w2419,w2418,w2417,w2416,w2415,w2414,w2413,w2412,w2411,w2410,w2409,w2408,w2407,w2406,w2405,w2404,w2403,w2402,w2401,w2400,w2399,w2398,w2397,w2396,w2395,w2394}, {w2614,w2613,w2612,w2611,w2610,w2609,w2608,w2607,w2606,w2605,w2604,w2603,w2602,w2601,w2600,w2599,w2598,w2597,w2596,w2595,w2594,w2593,w2592,w2591,w2590,w2589,w2588,w2587,w2586,w2585,w2584,w2583,w2582,w2581,w2580,w2579,w2578,w2577,w2576,w2575,w2574,w2573,w2572,w2571,w2570,w2569,w2568,w2567,w2566,w2565,w2564,w2563,w2562,w2561,w2560,w2559,w2558,w2557,w2556,w2555,w2554,w2553,w2552,w2551,w2550,w2549,w2548,w2547,w2546,w2545,w2544,w2543,w2542});
    wire w2905, w2906, w2907, w2908, w2978, w2979, w2980, w2981;
    sw_m #(.SIZE(73)) sw67({w2908,w2907,w2906,w2905,w2904,w2903,w2902,w2901,w2900,w2899,w2898,w2897,w2896,w2895,w2894,w2893,w2892,w2891,w2890,w2889,w2888,w2887,w2886,w2885,w2884,w2883,w2882,w2881,w2880,w2879,w2878,w2877,w2876,w2875,w2874,w2873,w2872,w2871,w2870,w2869,w2868,w2867,w2866,w2865,w2864,w2863,w2862,w2861,w2860,w2859,w2858,w2857,w2856,w2855,w2854,w2853,w2852,w2851,w2850,w2849,w2848,w2847,w2846,w2845,w2844,w2843,w2842,w2841,w2840,w2839,w2838,w2837,w2836}, {w2981,w2980,w2979,w2978,w2977,w2976,w2975,w2974,w2973,w2972,w2971,w2970,w2969,w2968,w2967,w2966,w2965,w2964,w2963,w2962,w2961,w2960,w2959,w2958,w2957,w2956,w2955,w2954,w2953,w2952,w2951,w2950,w2949,w2948,w2947,w2946,w2945,w2944,w2943,w2942,w2941,w2940,w2939,w2938,w2937,w2936,w2935,w2934,w2933,w2932,w2931,w2930,w2929,w2928,w2927,w2926,w2925,w2924,w2923,w2922,w2921,w2920,w2919,w2918,w2917,w2916,w2915,w2914,w2913,w2912,w2911,w2910,w2909}, w2541, {w2540,w2539,w2538,w2537,w2536,w2535,w2534,w2533,w2532,w2531,w2530,w2529,w2528,w2527,w2526,w2525,w2524,w2523,w2522,w2521,w2520,w2519,w2518,w2517,w2516,w2515,w2514,w2513,w2512,w2511,w2510,w2509,w2508,w2507,w2506,w2505,w2504,w2503,w2502,w2501,w2500,w2499,w2498,w2497,w2496,w2495,w2494,w2493,w2492,w2491,w2490,w2489,w2488,w2487,w2486,w2485,w2484,w2483,w2482,w2481,w2480,w2479,w2478,w2477,w2476,w2475,w2474,w2473,w2472,w2471,w2470,w2469,w2468}, {w2688,w2687,w2686,w2685,w2684,w2683,w2682,w2681,w2680,w2679,w2678,w2677,w2676,w2675,w2674,w2673,w2672,w2671,w2670,w2669,w2668,w2667,w2666,w2665,w2664,w2663,w2662,w2661,w2660,w2659,w2658,w2657,w2656,w2655,w2654,w2653,w2652,w2651,w2650,w2649,w2648,w2647,w2646,w2645,w2644,w2643,w2642,w2641,w2640,w2639,w2638,w2637,w2636,w2635,w2634,w2633,w2632,w2631,w2630,w2629,w2628,w2627,w2626,w2625,w2624,w2623,w2622,w2621,w2620,w2619,w2618,w2617,w2616});
    wire w3948, w3949, w3950, w3951, w4021, w4022, w4023, w4024;
    sw_m #(.SIZE(73)) sw68({w3951,w3950,w3949,w3948,w3947,w3946,w3945,w3944,w3943,w3942,w3941,w3940,w3939,w3938,w3937,w3936,w3935,w3934,w3933,w3932,w3931,w3930,w3929,w3928,w3927,w3926,w3925,w3924,w3923,w3922,w3921,w3920,w3919,w3918,w3917,w3916,w3915,w3914,w3913,w3912,w3911,w3910,w3909,w3908,w3907,w3906,w3905,w3904,w3903,w3902,w3901,w3900,w3899,w3898,w3897,w3896,w3895,w3894,w3893,w3892,w3891,w3890,w3889,w3888,w3887,w3886,w3885,w3884,w3883,w3882,w3881,w3880,w3879}, {w4024,w4023,w4022,w4021,w4020,w4019,w4018,w4017,w4016,w4015,w4014,w4013,w4012,w4011,w4010,w4009,w4008,w4007,w4006,w4005,w4004,w4003,w4002,w4001,w4000,w3999,w3998,w3997,w3996,w3995,w3994,w3993,w3992,w3991,w3990,w3989,w3988,w3987,w3986,w3985,w3984,w3983,w3982,w3981,w3980,w3979,w3978,w3977,w3976,w3975,w3974,w3973,w3972,w3971,w3970,w3969,w3968,w3967,w3966,w3965,w3964,w3963,w3962,w3961,w3960,w3959,w3958,w3957,w3956,w3955,w3954,w3953,w3952}, w3656, {w3655,w3654,w3653,w3652,w3651,w3650,w3649,w3648,w3647,w3646,w3645,w3644,w3643,w3642,w3641,w3640,w3639,w3638,w3637,w3636,w3635,w3634,w3633,w3632,w3631,w3630,w3629,w3628,w3627,w3626,w3625,w3624,w3623,w3622,w3621,w3620,w3619,w3618,w3617,w3616,w3615,w3614,w3613,w3612,w3611,w3610,w3609,w3608,w3607,w3606,w3605,w3604,w3603,w3602,w3601,w3600,w3599,w3598,w3597,w3596,w3595,w3594,w3593,w3592,w3591,w3590,w3589,w3588,w3587,w3586,w3585,w3584,w3583}, {w3803,w3802,w3801,w3800,w3799,w3798,w3797,w3796,w3795,w3794,w3793,w3792,w3791,w3790,w3789,w3788,w3787,w3786,w3785,w3784,w3783,w3782,w3781,w3780,w3779,w3778,w3777,w3776,w3775,w3774,w3773,w3772,w3771,w3770,w3769,w3768,w3767,w3766,w3765,w3764,w3763,w3762,w3761,w3760,w3759,w3758,w3757,w3756,w3755,w3754,w3753,w3752,w3751,w3750,w3749,w3748,w3747,w3746,w3745,w3744,w3743,w3742,w3741,w3740,w3739,w3738,w3737,w3736,w3735,w3734,w3733,w3732,w3731});
    wire w4094, w4095, w4096, w4097, w4167, w4168, w4169, w4170;
    sw_m #(.SIZE(73)) sw69({w4097,w4096,w4095,w4094,w4093,w4092,w4091,w4090,w4089,w4088,w4087,w4086,w4085,w4084,w4083,w4082,w4081,w4080,w4079,w4078,w4077,w4076,w4075,w4074,w4073,w4072,w4071,w4070,w4069,w4068,w4067,w4066,w4065,w4064,w4063,w4062,w4061,w4060,w4059,w4058,w4057,w4056,w4055,w4054,w4053,w4052,w4051,w4050,w4049,w4048,w4047,w4046,w4045,w4044,w4043,w4042,w4041,w4040,w4039,w4038,w4037,w4036,w4035,w4034,w4033,w4032,w4031,w4030,w4029,w4028,w4027,w4026,w4025}, {w4170,w4169,w4168,w4167,w4166,w4165,w4164,w4163,w4162,w4161,w4160,w4159,w4158,w4157,w4156,w4155,w4154,w4153,w4152,w4151,w4150,w4149,w4148,w4147,w4146,w4145,w4144,w4143,w4142,w4141,w4140,w4139,w4138,w4137,w4136,w4135,w4134,w4133,w4132,w4131,w4130,w4129,w4128,w4127,w4126,w4125,w4124,w4123,w4122,w4121,w4120,w4119,w4118,w4117,w4116,w4115,w4114,w4113,w4112,w4111,w4110,w4109,w4108,w4107,w4106,w4105,w4104,w4103,w4102,w4101,w4100,w4099,w4098}, w3730, {w3729,w3728,w3727,w3726,w3725,w3724,w3723,w3722,w3721,w3720,w3719,w3718,w3717,w3716,w3715,w3714,w3713,w3712,w3711,w3710,w3709,w3708,w3707,w3706,w3705,w3704,w3703,w3702,w3701,w3700,w3699,w3698,w3697,w3696,w3695,w3694,w3693,w3692,w3691,w3690,w3689,w3688,w3687,w3686,w3685,w3684,w3683,w3682,w3681,w3680,w3679,w3678,w3677,w3676,w3675,w3674,w3673,w3672,w3671,w3670,w3669,w3668,w3667,w3666,w3665,w3664,w3663,w3662,w3661,w3660,w3659,w3658,w3657}, {w3877,w3876,w3875,w3874,w3873,w3872,w3871,w3870,w3869,w3868,w3867,w3866,w3865,w3864,w3863,w3862,w3861,w3860,w3859,w3858,w3857,w3856,w3855,w3854,w3853,w3852,w3851,w3850,w3849,w3848,w3847,w3846,w3845,w3844,w3843,w3842,w3841,w3840,w3839,w3838,w3837,w3836,w3835,w3834,w3833,w3832,w3831,w3830,w3829,w3828,w3827,w3826,w3825,w3824,w3823,w3822,w3821,w3820,w3819,w3818,w3817,w3816,w3815,w3814,w3813,w3812,w3811,w3810,w3809,w3808,w3807,w3806,w3805});
    wire w4538, w4539, w4540, w4541, w4611, w4612, w4613, w4614;
    sw_m #(.SIZE(73)) sw70({w4541,w4540,w4539,w4538,w4537,w4536,w4535,w4534,w4533,w4532,w4531,w4530,w4529,w4528,w4527,w4526,w4525,w4524,w4523,w4522,w4521,w4520,w4519,w4518,w4517,w4516,w4515,w4514,w4513,w4512,w4511,w4510,w4509,w4508,w4507,w4506,w4505,w4504,w4503,w4502,w4501,w4500,w4499,w4498,w4497,w4496,w4495,w4494,w4493,w4492,w4491,w4490,w4489,w4488,w4487,w4486,w4485,w4484,w4483,w4482,w4481,w4480,w4479,w4478,w4477,w4476,w4475,w4474,w4473,w4472,w4471,w4470,w4469}, {w4614,w4613,w4612,w4611,w4610,w4609,w4608,w4607,w4606,w4605,w4604,w4603,w4602,w4601,w4600,w4599,w4598,w4597,w4596,w4595,w4594,w4593,w4592,w4591,w4590,w4589,w4588,w4587,w4586,w4585,w4584,w4583,w4582,w4581,w4580,w4579,w4578,w4577,w4576,w4575,w4574,w4573,w4572,w4571,w4570,w4569,w4568,w4567,w4566,w4565,w4564,w4563,w4562,w4561,w4560,w4559,w4558,w4557,w4556,w4555,w4554,w4553,w4552,w4551,w4550,w4549,w4548,w4547,w4546,w4545,w4544,w4543,w4542}, w4246, {w4245,w4244,w4243,w4242,w4241,w4240,w4239,w4238,w4237,w4236,w4235,w4234,w4233,w4232,w4231,w4230,w4229,w4228,w4227,w4226,w4225,w4224,w4223,w4222,w4221,w4220,w4219,w4218,w4217,w4216,w4215,w4214,w4213,w4212,w4211,w4210,w4209,w4208,w4207,w4206,w4205,w4204,w4203,w4202,w4201,w4200,w4199,w4198,w4197,w4196,w4195,w4194,w4193,w4192,w4191,w4190,w4189,w4188,w4187,w4186,w4185,w4184,w4183,w4182,w4181,w4180,w4179,w4178,w4177,w4176,w4175,w4174,w4173}, {w4393,w4392,w4391,w4390,w4389,w4388,w4387,w4386,w4385,w4384,w4383,w4382,w4381,w4380,w4379,w4378,w4377,w4376,w4375,w4374,w4373,w4372,w4371,w4370,w4369,w4368,w4367,w4366,w4365,w4364,w4363,w4362,w4361,w4360,w4359,w4358,w4357,w4356,w4355,w4354,w4353,w4352,w4351,w4350,w4349,w4348,w4347,w4346,w4345,w4344,w4343,w4342,w4341,w4340,w4339,w4338,w4337,w4336,w4335,w4334,w4333,w4332,w4331,w4330,w4329,w4328,w4327,w4326,w4325,w4324,w4323,w4322,w4321});
    wire w4684, w4685, w4686, w4687, w4757, w4758, w4759, w4760;
    sw_m #(.SIZE(73)) sw71({w4687,w4686,w4685,w4684,w4683,w4682,w4681,w4680,w4679,w4678,w4677,w4676,w4675,w4674,w4673,w4672,w4671,w4670,w4669,w4668,w4667,w4666,w4665,w4664,w4663,w4662,w4661,w4660,w4659,w4658,w4657,w4656,w4655,w4654,w4653,w4652,w4651,w4650,w4649,w4648,w4647,w4646,w4645,w4644,w4643,w4642,w4641,w4640,w4639,w4638,w4637,w4636,w4635,w4634,w4633,w4632,w4631,w4630,w4629,w4628,w4627,w4626,w4625,w4624,w4623,w4622,w4621,w4620,w4619,w4618,w4617,w4616,w4615}, {w4760,w4759,w4758,w4757,w4756,w4755,w4754,w4753,w4752,w4751,w4750,w4749,w4748,w4747,w4746,w4745,w4744,w4743,w4742,w4741,w4740,w4739,w4738,w4737,w4736,w4735,w4734,w4733,w4732,w4731,w4730,w4729,w4728,w4727,w4726,w4725,w4724,w4723,w4722,w4721,w4720,w4719,w4718,w4717,w4716,w4715,w4714,w4713,w4712,w4711,w4710,w4709,w4708,w4707,w4706,w4705,w4704,w4703,w4702,w4701,w4700,w4699,w4698,w4697,w4696,w4695,w4694,w4693,w4692,w4691,w4690,w4689,w4688}, w4320, {w4319,w4318,w4317,w4316,w4315,w4314,w4313,w4312,w4311,w4310,w4309,w4308,w4307,w4306,w4305,w4304,w4303,w4302,w4301,w4300,w4299,w4298,w4297,w4296,w4295,w4294,w4293,w4292,w4291,w4290,w4289,w4288,w4287,w4286,w4285,w4284,w4283,w4282,w4281,w4280,w4279,w4278,w4277,w4276,w4275,w4274,w4273,w4272,w4271,w4270,w4269,w4268,w4267,w4266,w4265,w4264,w4263,w4262,w4261,w4260,w4259,w4258,w4257,w4256,w4255,w4254,w4253,w4252,w4251,w4250,w4249,w4248,w4247}, {w4467,w4466,w4465,w4464,w4463,w4462,w4461,w4460,w4459,w4458,w4457,w4456,w4455,w4454,w4453,w4452,w4451,w4450,w4449,w4448,w4447,w4446,w4445,w4444,w4443,w4442,w4441,w4440,w4439,w4438,w4437,w4436,w4435,w4434,w4433,w4432,w4431,w4430,w4429,w4428,w4427,w4426,w4425,w4424,w4423,w4422,w4421,w4420,w4419,w4418,w4417,w4416,w4415,w4414,w4413,w4412,w4411,w4410,w4409,w4408,w4407,w4406,w4405,w4404,w4403,w4402,w4401,w4400,w4399,w4398,w4397,w4396,w4395});
    and and72(w4821, w2168, w2169);
    and and73(w4822, w2168, w2170);
    and and74(w4823, w2168, w2171);
    and and75(w4824, w2168, w2172);
    and and76(w4789, w2241, w2242);
    and and77(w4790, w2241, w2243);
    and and78(w4791, w2241, w2244);
    and and79(w4792, w2241, w2245);
    and and80(w4805, w2314, w2315);
    and and81(w4806, w2314, w2316);
    and and82(w4807, w2314, w2317);
    and and83(w4808, w2314, w2318);
    and and84(w4773, w2387, w2388);
    and and85(w4774, w2387, w2389);
    and and86(w4775, w2387, w2390);
    and and87(w4776, w2387, w2391);
    and and88(w4813, w2758, w2759);
    and and89(w4814, w2758, w2760);
    and and90(w4815, w2758, w2761);
    and and91(w4816, w2758, w2762);
    and and92(w4781, w2831, w2832);
    and and93(w4782, w2831, w2833);
    and and94(w4783, w2831, w2834);
    and and95(w4784, w2831, w2835);
    and and96(w4797, w2904, w2905);
    and and97(w4798, w2904, w2906);
    and and98(w4799, w2904, w2907);
    and and99(w4800, w2904, w2908);
    and and100(w4765, w2977, w2978);
    and and101(w4766, w2977, w2979);
    and and102(w4767, w2977, w2980);
    and and103(w4768, w2977, w2981);
    and and104(w4817, w3947, w3948);
    and and105(w4818, w3947, w3949);
    and and106(w4819, w3947, w3950);
    and and107(w4820, w3947, w3951);
    and and108(w4785, w4020, w4021);
    and and109(w4786, w4020, w4022);
    and and110(w4787, w4020, w4023);
    and and111(w4788, w4020, w4024);
    and and112(w4801, w4093, w4094);
    and and113(w4802, w4093, w4095);
    and and114(w4803, w4093, w4096);
    and and115(w4804, w4093, w4097);
    and and116(w4769, w4166, w4167);
    and and117(w4770, w4166, w4168);
    and and118(w4771, w4166, w4169);
    and and119(w4772, w4166, w4170);
    and and120(w4809, w4537, w4538);
    and and121(w4810, w4537, w4539);
    and and122(w4811, w4537, w4540);
    and and123(w4812, w4537, w4541);
    and and124(w4777, w4610, w4611);
    and and125(w4778, w4610, w4612);
    and and126(w4779, w4610, w4613);
    and and127(w4780, w4610, w4614);
    and and128(w4793, w4683, w4684);
    and and129(w4794, w4683, w4685);
    and and130(w4795, w4683, w4686);
    and and131(w4796, w4683, w4687);
    and and132(w4761, w4756, w4757);
    and and133(w4762, w4756, w4758);
    and and134(w4763, w4756, w4759);
    and and135(w4764, w4756, w4760);
endmodule
