`default_nettype none

module TNT_BIN_HC0_JaSJ17_68_16_4 (
output wire [69-1:0] out0,
output wire [69-1:0] out1,
output wire [69-1:0] out2,
output wire [69-1:0] out3,
output wire [69-1:0] out4,
output wire [69-1:0] out5,
output wire [69-1:0] out6,
output wire [69-1:0] out7,
output wire [69-1:0] out8,
output wire [69-1:0] out9,
output wire [69-1:0] out10,
output wire [69-1:0] out11,
output wire [69-1:0] out12,
output wire [69-1:0] out13,
output wire [69-1:0] out14,
output wire [69-1:0] out15,
input wire [70-1:0] in0,
input wire [70-1:0] in1,
input wire [70-1:0] in2,
input wire [70-1:0] in3,
input wire [70-1:0] in4,
input wire [70-1:0] in5,
input wire [70-1:0] in6,
input wire [70-1:0] in7,
input wire [70-1:0] in8,
input wire [70-1:0] in9,
input wire [70-1:0] in10,
input wire [70-1:0] in11,
input wire [70-1:0] in12,
input wire [70-1:0] in13,
input wire [70-1:0] in14,
input wire [70-1:0] in15);
    wire x0_0;
    wire x0_1;
    wire x0_2;
    wire x0_3;
    wire x0_4;
    wire x0_5;
    wire x0_6;
    wire x0_7;
    wire x0_8;
    wire x0_9;
    wire x0_10;
    wire x0_11;
    wire x0_12;
    wire x0_13;
    wire x0_14;
    wire x0_15;
    wire x0_16;
    wire x0_17;
    wire x0_18;
    wire x0_19;
    wire x0_20;
    wire x0_21;
    wire x0_22;
    wire x0_23;
    wire x0_24;
    wire x0_25;
    wire x0_26;
    wire x0_27;
    wire x0_28;
    wire x0_29;
    wire x0_30;
    wire x0_31;
    wire x0_32;
    wire x0_33;
    wire x0_34;
    wire x0_35;
    wire x0_36;
    wire x0_37;
    wire x0_38;
    wire x0_39;
    wire x0_40;
    wire x0_41;
    wire x0_42;
    wire x0_43;
    wire x0_44;
    wire x0_45;
    wire x0_46;
    wire x0_47;
    wire x0_48;
    wire x0_49;
    wire x0_50;
    wire x0_51;
    wire x0_52;
    wire x0_53;
    wire x0_54;
    wire x0_55;
    wire x0_56;
    wire x0_57;
    wire x0_58;
    wire x0_59;
    wire x0_60;
    wire x0_61;
    wire x0_62;
    wire x0_63;
    wire x0_64;
    wire x0_65;
    wire x0_66;
    wire x0_67;
    wire x0_68;
    wire x0_69;
    assign x0_0 = in0[0];
    assign x0_1 = in0[1];
    assign x0_2 = in0[2];
    assign x0_3 = in0[3];
    assign x0_4 = in0[4];
    assign x0_5 = in0[5];
    assign x0_6 = in0[6];
    assign x0_7 = in0[7];
    assign x0_8 = in0[8];
    assign x0_9 = in0[9];
    assign x0_10 = in0[10];
    assign x0_11 = in0[11];
    assign x0_12 = in0[12];
    assign x0_13 = in0[13];
    assign x0_14 = in0[14];
    assign x0_15 = in0[15];
    assign x0_16 = in0[16];
    assign x0_17 = in0[17];
    assign x0_18 = in0[18];
    assign x0_19 = in0[19];
    assign x0_20 = in0[20];
    assign x0_21 = in0[21];
    assign x0_22 = in0[22];
    assign x0_23 = in0[23];
    assign x0_24 = in0[24];
    assign x0_25 = in0[25];
    assign x0_26 = in0[26];
    assign x0_27 = in0[27];
    assign x0_28 = in0[28];
    assign x0_29 = in0[29];
    assign x0_30 = in0[30];
    assign x0_31 = in0[31];
    assign x0_32 = in0[32];
    assign x0_33 = in0[33];
    assign x0_34 = in0[34];
    assign x0_35 = in0[35];
    assign x0_36 = in0[36];
    assign x0_37 = in0[37];
    assign x0_38 = in0[38];
    assign x0_39 = in0[39];
    assign x0_40 = in0[40];
    assign x0_41 = in0[41];
    assign x0_42 = in0[42];
    assign x0_43 = in0[43];
    assign x0_44 = in0[44];
    assign x0_45 = in0[45];
    assign x0_46 = in0[46];
    assign x0_47 = in0[47];
    assign x0_48 = in0[48];
    assign x0_49 = in0[49];
    assign x0_50 = in0[50];
    assign x0_51 = in0[51];
    assign x0_52 = in0[52];
    assign x0_53 = in0[53];
    assign x0_54 = in0[54];
    assign x0_55 = in0[55];
    assign x0_56 = in0[56];
    assign x0_57 = in0[57];
    assign x0_58 = in0[58];
    assign x0_59 = in0[59];
    assign x0_60 = in0[60];
    assign x0_61 = in0[61];
    assign x0_62 = in0[62];
    assign x0_63 = in0[63];
    assign x0_64 = in0[64];
    assign x0_65 = in0[65];
    assign x0_66 = in0[66];
    assign x0_67 = in0[67];
    assign x0_68 = in0[68];
    assign x0_69 = in0[69];
    wire x1_0;
    wire x1_1;
    wire x1_2;
    wire x1_3;
    wire x1_4;
    wire x1_5;
    wire x1_6;
    wire x1_7;
    wire x1_8;
    wire x1_9;
    wire x1_10;
    wire x1_11;
    wire x1_12;
    wire x1_13;
    wire x1_14;
    wire x1_15;
    wire x1_16;
    wire x1_17;
    wire x1_18;
    wire x1_19;
    wire x1_20;
    wire x1_21;
    wire x1_22;
    wire x1_23;
    wire x1_24;
    wire x1_25;
    wire x1_26;
    wire x1_27;
    wire x1_28;
    wire x1_29;
    wire x1_30;
    wire x1_31;
    wire x1_32;
    wire x1_33;
    wire x1_34;
    wire x1_35;
    wire x1_36;
    wire x1_37;
    wire x1_38;
    wire x1_39;
    wire x1_40;
    wire x1_41;
    wire x1_42;
    wire x1_43;
    wire x1_44;
    wire x1_45;
    wire x1_46;
    wire x1_47;
    wire x1_48;
    wire x1_49;
    wire x1_50;
    wire x1_51;
    wire x1_52;
    wire x1_53;
    wire x1_54;
    wire x1_55;
    wire x1_56;
    wire x1_57;
    wire x1_58;
    wire x1_59;
    wire x1_60;
    wire x1_61;
    wire x1_62;
    wire x1_63;
    wire x1_64;
    wire x1_65;
    wire x1_66;
    wire x1_67;
    wire x1_68;
    wire x1_69;
    assign x1_0 = in1[0];
    assign x1_1 = in1[1];
    assign x1_2 = in1[2];
    assign x1_3 = in1[3];
    assign x1_4 = in1[4];
    assign x1_5 = in1[5];
    assign x1_6 = in1[6];
    assign x1_7 = in1[7];
    assign x1_8 = in1[8];
    assign x1_9 = in1[9];
    assign x1_10 = in1[10];
    assign x1_11 = in1[11];
    assign x1_12 = in1[12];
    assign x1_13 = in1[13];
    assign x1_14 = in1[14];
    assign x1_15 = in1[15];
    assign x1_16 = in1[16];
    assign x1_17 = in1[17];
    assign x1_18 = in1[18];
    assign x1_19 = in1[19];
    assign x1_20 = in1[20];
    assign x1_21 = in1[21];
    assign x1_22 = in1[22];
    assign x1_23 = in1[23];
    assign x1_24 = in1[24];
    assign x1_25 = in1[25];
    assign x1_26 = in1[26];
    assign x1_27 = in1[27];
    assign x1_28 = in1[28];
    assign x1_29 = in1[29];
    assign x1_30 = in1[30];
    assign x1_31 = in1[31];
    assign x1_32 = in1[32];
    assign x1_33 = in1[33];
    assign x1_34 = in1[34];
    assign x1_35 = in1[35];
    assign x1_36 = in1[36];
    assign x1_37 = in1[37];
    assign x1_38 = in1[38];
    assign x1_39 = in1[39];
    assign x1_40 = in1[40];
    assign x1_41 = in1[41];
    assign x1_42 = in1[42];
    assign x1_43 = in1[43];
    assign x1_44 = in1[44];
    assign x1_45 = in1[45];
    assign x1_46 = in1[46];
    assign x1_47 = in1[47];
    assign x1_48 = in1[48];
    assign x1_49 = in1[49];
    assign x1_50 = in1[50];
    assign x1_51 = in1[51];
    assign x1_52 = in1[52];
    assign x1_53 = in1[53];
    assign x1_54 = in1[54];
    assign x1_55 = in1[55];
    assign x1_56 = in1[56];
    assign x1_57 = in1[57];
    assign x1_58 = in1[58];
    assign x1_59 = in1[59];
    assign x1_60 = in1[60];
    assign x1_61 = in1[61];
    assign x1_62 = in1[62];
    assign x1_63 = in1[63];
    assign x1_64 = in1[64];
    assign x1_65 = in1[65];
    assign x1_66 = in1[66];
    assign x1_67 = in1[67];
    assign x1_68 = in1[68];
    assign x1_69 = in1[69];
    wire x2_0;
    wire x2_1;
    wire x2_2;
    wire x2_3;
    wire x2_4;
    wire x2_5;
    wire x2_6;
    wire x2_7;
    wire x2_8;
    wire x2_9;
    wire x2_10;
    wire x2_11;
    wire x2_12;
    wire x2_13;
    wire x2_14;
    wire x2_15;
    wire x2_16;
    wire x2_17;
    wire x2_18;
    wire x2_19;
    wire x2_20;
    wire x2_21;
    wire x2_22;
    wire x2_23;
    wire x2_24;
    wire x2_25;
    wire x2_26;
    wire x2_27;
    wire x2_28;
    wire x2_29;
    wire x2_30;
    wire x2_31;
    wire x2_32;
    wire x2_33;
    wire x2_34;
    wire x2_35;
    wire x2_36;
    wire x2_37;
    wire x2_38;
    wire x2_39;
    wire x2_40;
    wire x2_41;
    wire x2_42;
    wire x2_43;
    wire x2_44;
    wire x2_45;
    wire x2_46;
    wire x2_47;
    wire x2_48;
    wire x2_49;
    wire x2_50;
    wire x2_51;
    wire x2_52;
    wire x2_53;
    wire x2_54;
    wire x2_55;
    wire x2_56;
    wire x2_57;
    wire x2_58;
    wire x2_59;
    wire x2_60;
    wire x2_61;
    wire x2_62;
    wire x2_63;
    wire x2_64;
    wire x2_65;
    wire x2_66;
    wire x2_67;
    wire x2_68;
    wire x2_69;
    assign x2_0 = in2[0];
    assign x2_1 = in2[1];
    assign x2_2 = in2[2];
    assign x2_3 = in2[3];
    assign x2_4 = in2[4];
    assign x2_5 = in2[5];
    assign x2_6 = in2[6];
    assign x2_7 = in2[7];
    assign x2_8 = in2[8];
    assign x2_9 = in2[9];
    assign x2_10 = in2[10];
    assign x2_11 = in2[11];
    assign x2_12 = in2[12];
    assign x2_13 = in2[13];
    assign x2_14 = in2[14];
    assign x2_15 = in2[15];
    assign x2_16 = in2[16];
    assign x2_17 = in2[17];
    assign x2_18 = in2[18];
    assign x2_19 = in2[19];
    assign x2_20 = in2[20];
    assign x2_21 = in2[21];
    assign x2_22 = in2[22];
    assign x2_23 = in2[23];
    assign x2_24 = in2[24];
    assign x2_25 = in2[25];
    assign x2_26 = in2[26];
    assign x2_27 = in2[27];
    assign x2_28 = in2[28];
    assign x2_29 = in2[29];
    assign x2_30 = in2[30];
    assign x2_31 = in2[31];
    assign x2_32 = in2[32];
    assign x2_33 = in2[33];
    assign x2_34 = in2[34];
    assign x2_35 = in2[35];
    assign x2_36 = in2[36];
    assign x2_37 = in2[37];
    assign x2_38 = in2[38];
    assign x2_39 = in2[39];
    assign x2_40 = in2[40];
    assign x2_41 = in2[41];
    assign x2_42 = in2[42];
    assign x2_43 = in2[43];
    assign x2_44 = in2[44];
    assign x2_45 = in2[45];
    assign x2_46 = in2[46];
    assign x2_47 = in2[47];
    assign x2_48 = in2[48];
    assign x2_49 = in2[49];
    assign x2_50 = in2[50];
    assign x2_51 = in2[51];
    assign x2_52 = in2[52];
    assign x2_53 = in2[53];
    assign x2_54 = in2[54];
    assign x2_55 = in2[55];
    assign x2_56 = in2[56];
    assign x2_57 = in2[57];
    assign x2_58 = in2[58];
    assign x2_59 = in2[59];
    assign x2_60 = in2[60];
    assign x2_61 = in2[61];
    assign x2_62 = in2[62];
    assign x2_63 = in2[63];
    assign x2_64 = in2[64];
    assign x2_65 = in2[65];
    assign x2_66 = in2[66];
    assign x2_67 = in2[67];
    assign x2_68 = in2[68];
    assign x2_69 = in2[69];
    wire x3_0;
    wire x3_1;
    wire x3_2;
    wire x3_3;
    wire x3_4;
    wire x3_5;
    wire x3_6;
    wire x3_7;
    wire x3_8;
    wire x3_9;
    wire x3_10;
    wire x3_11;
    wire x3_12;
    wire x3_13;
    wire x3_14;
    wire x3_15;
    wire x3_16;
    wire x3_17;
    wire x3_18;
    wire x3_19;
    wire x3_20;
    wire x3_21;
    wire x3_22;
    wire x3_23;
    wire x3_24;
    wire x3_25;
    wire x3_26;
    wire x3_27;
    wire x3_28;
    wire x3_29;
    wire x3_30;
    wire x3_31;
    wire x3_32;
    wire x3_33;
    wire x3_34;
    wire x3_35;
    wire x3_36;
    wire x3_37;
    wire x3_38;
    wire x3_39;
    wire x3_40;
    wire x3_41;
    wire x3_42;
    wire x3_43;
    wire x3_44;
    wire x3_45;
    wire x3_46;
    wire x3_47;
    wire x3_48;
    wire x3_49;
    wire x3_50;
    wire x3_51;
    wire x3_52;
    wire x3_53;
    wire x3_54;
    wire x3_55;
    wire x3_56;
    wire x3_57;
    wire x3_58;
    wire x3_59;
    wire x3_60;
    wire x3_61;
    wire x3_62;
    wire x3_63;
    wire x3_64;
    wire x3_65;
    wire x3_66;
    wire x3_67;
    wire x3_68;
    wire x3_69;
    assign x3_0 = in3[0];
    assign x3_1 = in3[1];
    assign x3_2 = in3[2];
    assign x3_3 = in3[3];
    assign x3_4 = in3[4];
    assign x3_5 = in3[5];
    assign x3_6 = in3[6];
    assign x3_7 = in3[7];
    assign x3_8 = in3[8];
    assign x3_9 = in3[9];
    assign x3_10 = in3[10];
    assign x3_11 = in3[11];
    assign x3_12 = in3[12];
    assign x3_13 = in3[13];
    assign x3_14 = in3[14];
    assign x3_15 = in3[15];
    assign x3_16 = in3[16];
    assign x3_17 = in3[17];
    assign x3_18 = in3[18];
    assign x3_19 = in3[19];
    assign x3_20 = in3[20];
    assign x3_21 = in3[21];
    assign x3_22 = in3[22];
    assign x3_23 = in3[23];
    assign x3_24 = in3[24];
    assign x3_25 = in3[25];
    assign x3_26 = in3[26];
    assign x3_27 = in3[27];
    assign x3_28 = in3[28];
    assign x3_29 = in3[29];
    assign x3_30 = in3[30];
    assign x3_31 = in3[31];
    assign x3_32 = in3[32];
    assign x3_33 = in3[33];
    assign x3_34 = in3[34];
    assign x3_35 = in3[35];
    assign x3_36 = in3[36];
    assign x3_37 = in3[37];
    assign x3_38 = in3[38];
    assign x3_39 = in3[39];
    assign x3_40 = in3[40];
    assign x3_41 = in3[41];
    assign x3_42 = in3[42];
    assign x3_43 = in3[43];
    assign x3_44 = in3[44];
    assign x3_45 = in3[45];
    assign x3_46 = in3[46];
    assign x3_47 = in3[47];
    assign x3_48 = in3[48];
    assign x3_49 = in3[49];
    assign x3_50 = in3[50];
    assign x3_51 = in3[51];
    assign x3_52 = in3[52];
    assign x3_53 = in3[53];
    assign x3_54 = in3[54];
    assign x3_55 = in3[55];
    assign x3_56 = in3[56];
    assign x3_57 = in3[57];
    assign x3_58 = in3[58];
    assign x3_59 = in3[59];
    assign x3_60 = in3[60];
    assign x3_61 = in3[61];
    assign x3_62 = in3[62];
    assign x3_63 = in3[63];
    assign x3_64 = in3[64];
    assign x3_65 = in3[65];
    assign x3_66 = in3[66];
    assign x3_67 = in3[67];
    assign x3_68 = in3[68];
    assign x3_69 = in3[69];
    wire x4_0;
    wire x4_1;
    wire x4_2;
    wire x4_3;
    wire x4_4;
    wire x4_5;
    wire x4_6;
    wire x4_7;
    wire x4_8;
    wire x4_9;
    wire x4_10;
    wire x4_11;
    wire x4_12;
    wire x4_13;
    wire x4_14;
    wire x4_15;
    wire x4_16;
    wire x4_17;
    wire x4_18;
    wire x4_19;
    wire x4_20;
    wire x4_21;
    wire x4_22;
    wire x4_23;
    wire x4_24;
    wire x4_25;
    wire x4_26;
    wire x4_27;
    wire x4_28;
    wire x4_29;
    wire x4_30;
    wire x4_31;
    wire x4_32;
    wire x4_33;
    wire x4_34;
    wire x4_35;
    wire x4_36;
    wire x4_37;
    wire x4_38;
    wire x4_39;
    wire x4_40;
    wire x4_41;
    wire x4_42;
    wire x4_43;
    wire x4_44;
    wire x4_45;
    wire x4_46;
    wire x4_47;
    wire x4_48;
    wire x4_49;
    wire x4_50;
    wire x4_51;
    wire x4_52;
    wire x4_53;
    wire x4_54;
    wire x4_55;
    wire x4_56;
    wire x4_57;
    wire x4_58;
    wire x4_59;
    wire x4_60;
    wire x4_61;
    wire x4_62;
    wire x4_63;
    wire x4_64;
    wire x4_65;
    wire x4_66;
    wire x4_67;
    wire x4_68;
    wire x4_69;
    assign x4_0 = in4[0];
    assign x4_1 = in4[1];
    assign x4_2 = in4[2];
    assign x4_3 = in4[3];
    assign x4_4 = in4[4];
    assign x4_5 = in4[5];
    assign x4_6 = in4[6];
    assign x4_7 = in4[7];
    assign x4_8 = in4[8];
    assign x4_9 = in4[9];
    assign x4_10 = in4[10];
    assign x4_11 = in4[11];
    assign x4_12 = in4[12];
    assign x4_13 = in4[13];
    assign x4_14 = in4[14];
    assign x4_15 = in4[15];
    assign x4_16 = in4[16];
    assign x4_17 = in4[17];
    assign x4_18 = in4[18];
    assign x4_19 = in4[19];
    assign x4_20 = in4[20];
    assign x4_21 = in4[21];
    assign x4_22 = in4[22];
    assign x4_23 = in4[23];
    assign x4_24 = in4[24];
    assign x4_25 = in4[25];
    assign x4_26 = in4[26];
    assign x4_27 = in4[27];
    assign x4_28 = in4[28];
    assign x4_29 = in4[29];
    assign x4_30 = in4[30];
    assign x4_31 = in4[31];
    assign x4_32 = in4[32];
    assign x4_33 = in4[33];
    assign x4_34 = in4[34];
    assign x4_35 = in4[35];
    assign x4_36 = in4[36];
    assign x4_37 = in4[37];
    assign x4_38 = in4[38];
    assign x4_39 = in4[39];
    assign x4_40 = in4[40];
    assign x4_41 = in4[41];
    assign x4_42 = in4[42];
    assign x4_43 = in4[43];
    assign x4_44 = in4[44];
    assign x4_45 = in4[45];
    assign x4_46 = in4[46];
    assign x4_47 = in4[47];
    assign x4_48 = in4[48];
    assign x4_49 = in4[49];
    assign x4_50 = in4[50];
    assign x4_51 = in4[51];
    assign x4_52 = in4[52];
    assign x4_53 = in4[53];
    assign x4_54 = in4[54];
    assign x4_55 = in4[55];
    assign x4_56 = in4[56];
    assign x4_57 = in4[57];
    assign x4_58 = in4[58];
    assign x4_59 = in4[59];
    assign x4_60 = in4[60];
    assign x4_61 = in4[61];
    assign x4_62 = in4[62];
    assign x4_63 = in4[63];
    assign x4_64 = in4[64];
    assign x4_65 = in4[65];
    assign x4_66 = in4[66];
    assign x4_67 = in4[67];
    assign x4_68 = in4[68];
    assign x4_69 = in4[69];
    wire x5_0;
    wire x5_1;
    wire x5_2;
    wire x5_3;
    wire x5_4;
    wire x5_5;
    wire x5_6;
    wire x5_7;
    wire x5_8;
    wire x5_9;
    wire x5_10;
    wire x5_11;
    wire x5_12;
    wire x5_13;
    wire x5_14;
    wire x5_15;
    wire x5_16;
    wire x5_17;
    wire x5_18;
    wire x5_19;
    wire x5_20;
    wire x5_21;
    wire x5_22;
    wire x5_23;
    wire x5_24;
    wire x5_25;
    wire x5_26;
    wire x5_27;
    wire x5_28;
    wire x5_29;
    wire x5_30;
    wire x5_31;
    wire x5_32;
    wire x5_33;
    wire x5_34;
    wire x5_35;
    wire x5_36;
    wire x5_37;
    wire x5_38;
    wire x5_39;
    wire x5_40;
    wire x5_41;
    wire x5_42;
    wire x5_43;
    wire x5_44;
    wire x5_45;
    wire x5_46;
    wire x5_47;
    wire x5_48;
    wire x5_49;
    wire x5_50;
    wire x5_51;
    wire x5_52;
    wire x5_53;
    wire x5_54;
    wire x5_55;
    wire x5_56;
    wire x5_57;
    wire x5_58;
    wire x5_59;
    wire x5_60;
    wire x5_61;
    wire x5_62;
    wire x5_63;
    wire x5_64;
    wire x5_65;
    wire x5_66;
    wire x5_67;
    wire x5_68;
    wire x5_69;
    assign x5_0 = in5[0];
    assign x5_1 = in5[1];
    assign x5_2 = in5[2];
    assign x5_3 = in5[3];
    assign x5_4 = in5[4];
    assign x5_5 = in5[5];
    assign x5_6 = in5[6];
    assign x5_7 = in5[7];
    assign x5_8 = in5[8];
    assign x5_9 = in5[9];
    assign x5_10 = in5[10];
    assign x5_11 = in5[11];
    assign x5_12 = in5[12];
    assign x5_13 = in5[13];
    assign x5_14 = in5[14];
    assign x5_15 = in5[15];
    assign x5_16 = in5[16];
    assign x5_17 = in5[17];
    assign x5_18 = in5[18];
    assign x5_19 = in5[19];
    assign x5_20 = in5[20];
    assign x5_21 = in5[21];
    assign x5_22 = in5[22];
    assign x5_23 = in5[23];
    assign x5_24 = in5[24];
    assign x5_25 = in5[25];
    assign x5_26 = in5[26];
    assign x5_27 = in5[27];
    assign x5_28 = in5[28];
    assign x5_29 = in5[29];
    assign x5_30 = in5[30];
    assign x5_31 = in5[31];
    assign x5_32 = in5[32];
    assign x5_33 = in5[33];
    assign x5_34 = in5[34];
    assign x5_35 = in5[35];
    assign x5_36 = in5[36];
    assign x5_37 = in5[37];
    assign x5_38 = in5[38];
    assign x5_39 = in5[39];
    assign x5_40 = in5[40];
    assign x5_41 = in5[41];
    assign x5_42 = in5[42];
    assign x5_43 = in5[43];
    assign x5_44 = in5[44];
    assign x5_45 = in5[45];
    assign x5_46 = in5[46];
    assign x5_47 = in5[47];
    assign x5_48 = in5[48];
    assign x5_49 = in5[49];
    assign x5_50 = in5[50];
    assign x5_51 = in5[51];
    assign x5_52 = in5[52];
    assign x5_53 = in5[53];
    assign x5_54 = in5[54];
    assign x5_55 = in5[55];
    assign x5_56 = in5[56];
    assign x5_57 = in5[57];
    assign x5_58 = in5[58];
    assign x5_59 = in5[59];
    assign x5_60 = in5[60];
    assign x5_61 = in5[61];
    assign x5_62 = in5[62];
    assign x5_63 = in5[63];
    assign x5_64 = in5[64];
    assign x5_65 = in5[65];
    assign x5_66 = in5[66];
    assign x5_67 = in5[67];
    assign x5_68 = in5[68];
    assign x5_69 = in5[69];
    wire x6_0;
    wire x6_1;
    wire x6_2;
    wire x6_3;
    wire x6_4;
    wire x6_5;
    wire x6_6;
    wire x6_7;
    wire x6_8;
    wire x6_9;
    wire x6_10;
    wire x6_11;
    wire x6_12;
    wire x6_13;
    wire x6_14;
    wire x6_15;
    wire x6_16;
    wire x6_17;
    wire x6_18;
    wire x6_19;
    wire x6_20;
    wire x6_21;
    wire x6_22;
    wire x6_23;
    wire x6_24;
    wire x6_25;
    wire x6_26;
    wire x6_27;
    wire x6_28;
    wire x6_29;
    wire x6_30;
    wire x6_31;
    wire x6_32;
    wire x6_33;
    wire x6_34;
    wire x6_35;
    wire x6_36;
    wire x6_37;
    wire x6_38;
    wire x6_39;
    wire x6_40;
    wire x6_41;
    wire x6_42;
    wire x6_43;
    wire x6_44;
    wire x6_45;
    wire x6_46;
    wire x6_47;
    wire x6_48;
    wire x6_49;
    wire x6_50;
    wire x6_51;
    wire x6_52;
    wire x6_53;
    wire x6_54;
    wire x6_55;
    wire x6_56;
    wire x6_57;
    wire x6_58;
    wire x6_59;
    wire x6_60;
    wire x6_61;
    wire x6_62;
    wire x6_63;
    wire x6_64;
    wire x6_65;
    wire x6_66;
    wire x6_67;
    wire x6_68;
    wire x6_69;
    assign x6_0 = in6[0];
    assign x6_1 = in6[1];
    assign x6_2 = in6[2];
    assign x6_3 = in6[3];
    assign x6_4 = in6[4];
    assign x6_5 = in6[5];
    assign x6_6 = in6[6];
    assign x6_7 = in6[7];
    assign x6_8 = in6[8];
    assign x6_9 = in6[9];
    assign x6_10 = in6[10];
    assign x6_11 = in6[11];
    assign x6_12 = in6[12];
    assign x6_13 = in6[13];
    assign x6_14 = in6[14];
    assign x6_15 = in6[15];
    assign x6_16 = in6[16];
    assign x6_17 = in6[17];
    assign x6_18 = in6[18];
    assign x6_19 = in6[19];
    assign x6_20 = in6[20];
    assign x6_21 = in6[21];
    assign x6_22 = in6[22];
    assign x6_23 = in6[23];
    assign x6_24 = in6[24];
    assign x6_25 = in6[25];
    assign x6_26 = in6[26];
    assign x6_27 = in6[27];
    assign x6_28 = in6[28];
    assign x6_29 = in6[29];
    assign x6_30 = in6[30];
    assign x6_31 = in6[31];
    assign x6_32 = in6[32];
    assign x6_33 = in6[33];
    assign x6_34 = in6[34];
    assign x6_35 = in6[35];
    assign x6_36 = in6[36];
    assign x6_37 = in6[37];
    assign x6_38 = in6[38];
    assign x6_39 = in6[39];
    assign x6_40 = in6[40];
    assign x6_41 = in6[41];
    assign x6_42 = in6[42];
    assign x6_43 = in6[43];
    assign x6_44 = in6[44];
    assign x6_45 = in6[45];
    assign x6_46 = in6[46];
    assign x6_47 = in6[47];
    assign x6_48 = in6[48];
    assign x6_49 = in6[49];
    assign x6_50 = in6[50];
    assign x6_51 = in6[51];
    assign x6_52 = in6[52];
    assign x6_53 = in6[53];
    assign x6_54 = in6[54];
    assign x6_55 = in6[55];
    assign x6_56 = in6[56];
    assign x6_57 = in6[57];
    assign x6_58 = in6[58];
    assign x6_59 = in6[59];
    assign x6_60 = in6[60];
    assign x6_61 = in6[61];
    assign x6_62 = in6[62];
    assign x6_63 = in6[63];
    assign x6_64 = in6[64];
    assign x6_65 = in6[65];
    assign x6_66 = in6[66];
    assign x6_67 = in6[67];
    assign x6_68 = in6[68];
    assign x6_69 = in6[69];
    wire x7_0;
    wire x7_1;
    wire x7_2;
    wire x7_3;
    wire x7_4;
    wire x7_5;
    wire x7_6;
    wire x7_7;
    wire x7_8;
    wire x7_9;
    wire x7_10;
    wire x7_11;
    wire x7_12;
    wire x7_13;
    wire x7_14;
    wire x7_15;
    wire x7_16;
    wire x7_17;
    wire x7_18;
    wire x7_19;
    wire x7_20;
    wire x7_21;
    wire x7_22;
    wire x7_23;
    wire x7_24;
    wire x7_25;
    wire x7_26;
    wire x7_27;
    wire x7_28;
    wire x7_29;
    wire x7_30;
    wire x7_31;
    wire x7_32;
    wire x7_33;
    wire x7_34;
    wire x7_35;
    wire x7_36;
    wire x7_37;
    wire x7_38;
    wire x7_39;
    wire x7_40;
    wire x7_41;
    wire x7_42;
    wire x7_43;
    wire x7_44;
    wire x7_45;
    wire x7_46;
    wire x7_47;
    wire x7_48;
    wire x7_49;
    wire x7_50;
    wire x7_51;
    wire x7_52;
    wire x7_53;
    wire x7_54;
    wire x7_55;
    wire x7_56;
    wire x7_57;
    wire x7_58;
    wire x7_59;
    wire x7_60;
    wire x7_61;
    wire x7_62;
    wire x7_63;
    wire x7_64;
    wire x7_65;
    wire x7_66;
    wire x7_67;
    wire x7_68;
    wire x7_69;
    assign x7_0 = in7[0];
    assign x7_1 = in7[1];
    assign x7_2 = in7[2];
    assign x7_3 = in7[3];
    assign x7_4 = in7[4];
    assign x7_5 = in7[5];
    assign x7_6 = in7[6];
    assign x7_7 = in7[7];
    assign x7_8 = in7[8];
    assign x7_9 = in7[9];
    assign x7_10 = in7[10];
    assign x7_11 = in7[11];
    assign x7_12 = in7[12];
    assign x7_13 = in7[13];
    assign x7_14 = in7[14];
    assign x7_15 = in7[15];
    assign x7_16 = in7[16];
    assign x7_17 = in7[17];
    assign x7_18 = in7[18];
    assign x7_19 = in7[19];
    assign x7_20 = in7[20];
    assign x7_21 = in7[21];
    assign x7_22 = in7[22];
    assign x7_23 = in7[23];
    assign x7_24 = in7[24];
    assign x7_25 = in7[25];
    assign x7_26 = in7[26];
    assign x7_27 = in7[27];
    assign x7_28 = in7[28];
    assign x7_29 = in7[29];
    assign x7_30 = in7[30];
    assign x7_31 = in7[31];
    assign x7_32 = in7[32];
    assign x7_33 = in7[33];
    assign x7_34 = in7[34];
    assign x7_35 = in7[35];
    assign x7_36 = in7[36];
    assign x7_37 = in7[37];
    assign x7_38 = in7[38];
    assign x7_39 = in7[39];
    assign x7_40 = in7[40];
    assign x7_41 = in7[41];
    assign x7_42 = in7[42];
    assign x7_43 = in7[43];
    assign x7_44 = in7[44];
    assign x7_45 = in7[45];
    assign x7_46 = in7[46];
    assign x7_47 = in7[47];
    assign x7_48 = in7[48];
    assign x7_49 = in7[49];
    assign x7_50 = in7[50];
    assign x7_51 = in7[51];
    assign x7_52 = in7[52];
    assign x7_53 = in7[53];
    assign x7_54 = in7[54];
    assign x7_55 = in7[55];
    assign x7_56 = in7[56];
    assign x7_57 = in7[57];
    assign x7_58 = in7[58];
    assign x7_59 = in7[59];
    assign x7_60 = in7[60];
    assign x7_61 = in7[61];
    assign x7_62 = in7[62];
    assign x7_63 = in7[63];
    assign x7_64 = in7[64];
    assign x7_65 = in7[65];
    assign x7_66 = in7[66];
    assign x7_67 = in7[67];
    assign x7_68 = in7[68];
    assign x7_69 = in7[69];
    wire x8_0;
    wire x8_1;
    wire x8_2;
    wire x8_3;
    wire x8_4;
    wire x8_5;
    wire x8_6;
    wire x8_7;
    wire x8_8;
    wire x8_9;
    wire x8_10;
    wire x8_11;
    wire x8_12;
    wire x8_13;
    wire x8_14;
    wire x8_15;
    wire x8_16;
    wire x8_17;
    wire x8_18;
    wire x8_19;
    wire x8_20;
    wire x8_21;
    wire x8_22;
    wire x8_23;
    wire x8_24;
    wire x8_25;
    wire x8_26;
    wire x8_27;
    wire x8_28;
    wire x8_29;
    wire x8_30;
    wire x8_31;
    wire x8_32;
    wire x8_33;
    wire x8_34;
    wire x8_35;
    wire x8_36;
    wire x8_37;
    wire x8_38;
    wire x8_39;
    wire x8_40;
    wire x8_41;
    wire x8_42;
    wire x8_43;
    wire x8_44;
    wire x8_45;
    wire x8_46;
    wire x8_47;
    wire x8_48;
    wire x8_49;
    wire x8_50;
    wire x8_51;
    wire x8_52;
    wire x8_53;
    wire x8_54;
    wire x8_55;
    wire x8_56;
    wire x8_57;
    wire x8_58;
    wire x8_59;
    wire x8_60;
    wire x8_61;
    wire x8_62;
    wire x8_63;
    wire x8_64;
    wire x8_65;
    wire x8_66;
    wire x8_67;
    wire x8_68;
    wire x8_69;
    assign x8_0 = in8[0];
    assign x8_1 = in8[1];
    assign x8_2 = in8[2];
    assign x8_3 = in8[3];
    assign x8_4 = in8[4];
    assign x8_5 = in8[5];
    assign x8_6 = in8[6];
    assign x8_7 = in8[7];
    assign x8_8 = in8[8];
    assign x8_9 = in8[9];
    assign x8_10 = in8[10];
    assign x8_11 = in8[11];
    assign x8_12 = in8[12];
    assign x8_13 = in8[13];
    assign x8_14 = in8[14];
    assign x8_15 = in8[15];
    assign x8_16 = in8[16];
    assign x8_17 = in8[17];
    assign x8_18 = in8[18];
    assign x8_19 = in8[19];
    assign x8_20 = in8[20];
    assign x8_21 = in8[21];
    assign x8_22 = in8[22];
    assign x8_23 = in8[23];
    assign x8_24 = in8[24];
    assign x8_25 = in8[25];
    assign x8_26 = in8[26];
    assign x8_27 = in8[27];
    assign x8_28 = in8[28];
    assign x8_29 = in8[29];
    assign x8_30 = in8[30];
    assign x8_31 = in8[31];
    assign x8_32 = in8[32];
    assign x8_33 = in8[33];
    assign x8_34 = in8[34];
    assign x8_35 = in8[35];
    assign x8_36 = in8[36];
    assign x8_37 = in8[37];
    assign x8_38 = in8[38];
    assign x8_39 = in8[39];
    assign x8_40 = in8[40];
    assign x8_41 = in8[41];
    assign x8_42 = in8[42];
    assign x8_43 = in8[43];
    assign x8_44 = in8[44];
    assign x8_45 = in8[45];
    assign x8_46 = in8[46];
    assign x8_47 = in8[47];
    assign x8_48 = in8[48];
    assign x8_49 = in8[49];
    assign x8_50 = in8[50];
    assign x8_51 = in8[51];
    assign x8_52 = in8[52];
    assign x8_53 = in8[53];
    assign x8_54 = in8[54];
    assign x8_55 = in8[55];
    assign x8_56 = in8[56];
    assign x8_57 = in8[57];
    assign x8_58 = in8[58];
    assign x8_59 = in8[59];
    assign x8_60 = in8[60];
    assign x8_61 = in8[61];
    assign x8_62 = in8[62];
    assign x8_63 = in8[63];
    assign x8_64 = in8[64];
    assign x8_65 = in8[65];
    assign x8_66 = in8[66];
    assign x8_67 = in8[67];
    assign x8_68 = in8[68];
    assign x8_69 = in8[69];
    wire x9_0;
    wire x9_1;
    wire x9_2;
    wire x9_3;
    wire x9_4;
    wire x9_5;
    wire x9_6;
    wire x9_7;
    wire x9_8;
    wire x9_9;
    wire x9_10;
    wire x9_11;
    wire x9_12;
    wire x9_13;
    wire x9_14;
    wire x9_15;
    wire x9_16;
    wire x9_17;
    wire x9_18;
    wire x9_19;
    wire x9_20;
    wire x9_21;
    wire x9_22;
    wire x9_23;
    wire x9_24;
    wire x9_25;
    wire x9_26;
    wire x9_27;
    wire x9_28;
    wire x9_29;
    wire x9_30;
    wire x9_31;
    wire x9_32;
    wire x9_33;
    wire x9_34;
    wire x9_35;
    wire x9_36;
    wire x9_37;
    wire x9_38;
    wire x9_39;
    wire x9_40;
    wire x9_41;
    wire x9_42;
    wire x9_43;
    wire x9_44;
    wire x9_45;
    wire x9_46;
    wire x9_47;
    wire x9_48;
    wire x9_49;
    wire x9_50;
    wire x9_51;
    wire x9_52;
    wire x9_53;
    wire x9_54;
    wire x9_55;
    wire x9_56;
    wire x9_57;
    wire x9_58;
    wire x9_59;
    wire x9_60;
    wire x9_61;
    wire x9_62;
    wire x9_63;
    wire x9_64;
    wire x9_65;
    wire x9_66;
    wire x9_67;
    wire x9_68;
    wire x9_69;
    assign x9_0 = in9[0];
    assign x9_1 = in9[1];
    assign x9_2 = in9[2];
    assign x9_3 = in9[3];
    assign x9_4 = in9[4];
    assign x9_5 = in9[5];
    assign x9_6 = in9[6];
    assign x9_7 = in9[7];
    assign x9_8 = in9[8];
    assign x9_9 = in9[9];
    assign x9_10 = in9[10];
    assign x9_11 = in9[11];
    assign x9_12 = in9[12];
    assign x9_13 = in9[13];
    assign x9_14 = in9[14];
    assign x9_15 = in9[15];
    assign x9_16 = in9[16];
    assign x9_17 = in9[17];
    assign x9_18 = in9[18];
    assign x9_19 = in9[19];
    assign x9_20 = in9[20];
    assign x9_21 = in9[21];
    assign x9_22 = in9[22];
    assign x9_23 = in9[23];
    assign x9_24 = in9[24];
    assign x9_25 = in9[25];
    assign x9_26 = in9[26];
    assign x9_27 = in9[27];
    assign x9_28 = in9[28];
    assign x9_29 = in9[29];
    assign x9_30 = in9[30];
    assign x9_31 = in9[31];
    assign x9_32 = in9[32];
    assign x9_33 = in9[33];
    assign x9_34 = in9[34];
    assign x9_35 = in9[35];
    assign x9_36 = in9[36];
    assign x9_37 = in9[37];
    assign x9_38 = in9[38];
    assign x9_39 = in9[39];
    assign x9_40 = in9[40];
    assign x9_41 = in9[41];
    assign x9_42 = in9[42];
    assign x9_43 = in9[43];
    assign x9_44 = in9[44];
    assign x9_45 = in9[45];
    assign x9_46 = in9[46];
    assign x9_47 = in9[47];
    assign x9_48 = in9[48];
    assign x9_49 = in9[49];
    assign x9_50 = in9[50];
    assign x9_51 = in9[51];
    assign x9_52 = in9[52];
    assign x9_53 = in9[53];
    assign x9_54 = in9[54];
    assign x9_55 = in9[55];
    assign x9_56 = in9[56];
    assign x9_57 = in9[57];
    assign x9_58 = in9[58];
    assign x9_59 = in9[59];
    assign x9_60 = in9[60];
    assign x9_61 = in9[61];
    assign x9_62 = in9[62];
    assign x9_63 = in9[63];
    assign x9_64 = in9[64];
    assign x9_65 = in9[65];
    assign x9_66 = in9[66];
    assign x9_67 = in9[67];
    assign x9_68 = in9[68];
    assign x9_69 = in9[69];
    wire x10_0;
    wire x10_1;
    wire x10_2;
    wire x10_3;
    wire x10_4;
    wire x10_5;
    wire x10_6;
    wire x10_7;
    wire x10_8;
    wire x10_9;
    wire x10_10;
    wire x10_11;
    wire x10_12;
    wire x10_13;
    wire x10_14;
    wire x10_15;
    wire x10_16;
    wire x10_17;
    wire x10_18;
    wire x10_19;
    wire x10_20;
    wire x10_21;
    wire x10_22;
    wire x10_23;
    wire x10_24;
    wire x10_25;
    wire x10_26;
    wire x10_27;
    wire x10_28;
    wire x10_29;
    wire x10_30;
    wire x10_31;
    wire x10_32;
    wire x10_33;
    wire x10_34;
    wire x10_35;
    wire x10_36;
    wire x10_37;
    wire x10_38;
    wire x10_39;
    wire x10_40;
    wire x10_41;
    wire x10_42;
    wire x10_43;
    wire x10_44;
    wire x10_45;
    wire x10_46;
    wire x10_47;
    wire x10_48;
    wire x10_49;
    wire x10_50;
    wire x10_51;
    wire x10_52;
    wire x10_53;
    wire x10_54;
    wire x10_55;
    wire x10_56;
    wire x10_57;
    wire x10_58;
    wire x10_59;
    wire x10_60;
    wire x10_61;
    wire x10_62;
    wire x10_63;
    wire x10_64;
    wire x10_65;
    wire x10_66;
    wire x10_67;
    wire x10_68;
    wire x10_69;
    assign x10_0 = in10[0];
    assign x10_1 = in10[1];
    assign x10_2 = in10[2];
    assign x10_3 = in10[3];
    assign x10_4 = in10[4];
    assign x10_5 = in10[5];
    assign x10_6 = in10[6];
    assign x10_7 = in10[7];
    assign x10_8 = in10[8];
    assign x10_9 = in10[9];
    assign x10_10 = in10[10];
    assign x10_11 = in10[11];
    assign x10_12 = in10[12];
    assign x10_13 = in10[13];
    assign x10_14 = in10[14];
    assign x10_15 = in10[15];
    assign x10_16 = in10[16];
    assign x10_17 = in10[17];
    assign x10_18 = in10[18];
    assign x10_19 = in10[19];
    assign x10_20 = in10[20];
    assign x10_21 = in10[21];
    assign x10_22 = in10[22];
    assign x10_23 = in10[23];
    assign x10_24 = in10[24];
    assign x10_25 = in10[25];
    assign x10_26 = in10[26];
    assign x10_27 = in10[27];
    assign x10_28 = in10[28];
    assign x10_29 = in10[29];
    assign x10_30 = in10[30];
    assign x10_31 = in10[31];
    assign x10_32 = in10[32];
    assign x10_33 = in10[33];
    assign x10_34 = in10[34];
    assign x10_35 = in10[35];
    assign x10_36 = in10[36];
    assign x10_37 = in10[37];
    assign x10_38 = in10[38];
    assign x10_39 = in10[39];
    assign x10_40 = in10[40];
    assign x10_41 = in10[41];
    assign x10_42 = in10[42];
    assign x10_43 = in10[43];
    assign x10_44 = in10[44];
    assign x10_45 = in10[45];
    assign x10_46 = in10[46];
    assign x10_47 = in10[47];
    assign x10_48 = in10[48];
    assign x10_49 = in10[49];
    assign x10_50 = in10[50];
    assign x10_51 = in10[51];
    assign x10_52 = in10[52];
    assign x10_53 = in10[53];
    assign x10_54 = in10[54];
    assign x10_55 = in10[55];
    assign x10_56 = in10[56];
    assign x10_57 = in10[57];
    assign x10_58 = in10[58];
    assign x10_59 = in10[59];
    assign x10_60 = in10[60];
    assign x10_61 = in10[61];
    assign x10_62 = in10[62];
    assign x10_63 = in10[63];
    assign x10_64 = in10[64];
    assign x10_65 = in10[65];
    assign x10_66 = in10[66];
    assign x10_67 = in10[67];
    assign x10_68 = in10[68];
    assign x10_69 = in10[69];
    wire x11_0;
    wire x11_1;
    wire x11_2;
    wire x11_3;
    wire x11_4;
    wire x11_5;
    wire x11_6;
    wire x11_7;
    wire x11_8;
    wire x11_9;
    wire x11_10;
    wire x11_11;
    wire x11_12;
    wire x11_13;
    wire x11_14;
    wire x11_15;
    wire x11_16;
    wire x11_17;
    wire x11_18;
    wire x11_19;
    wire x11_20;
    wire x11_21;
    wire x11_22;
    wire x11_23;
    wire x11_24;
    wire x11_25;
    wire x11_26;
    wire x11_27;
    wire x11_28;
    wire x11_29;
    wire x11_30;
    wire x11_31;
    wire x11_32;
    wire x11_33;
    wire x11_34;
    wire x11_35;
    wire x11_36;
    wire x11_37;
    wire x11_38;
    wire x11_39;
    wire x11_40;
    wire x11_41;
    wire x11_42;
    wire x11_43;
    wire x11_44;
    wire x11_45;
    wire x11_46;
    wire x11_47;
    wire x11_48;
    wire x11_49;
    wire x11_50;
    wire x11_51;
    wire x11_52;
    wire x11_53;
    wire x11_54;
    wire x11_55;
    wire x11_56;
    wire x11_57;
    wire x11_58;
    wire x11_59;
    wire x11_60;
    wire x11_61;
    wire x11_62;
    wire x11_63;
    wire x11_64;
    wire x11_65;
    wire x11_66;
    wire x11_67;
    wire x11_68;
    wire x11_69;
    assign x11_0 = in11[0];
    assign x11_1 = in11[1];
    assign x11_2 = in11[2];
    assign x11_3 = in11[3];
    assign x11_4 = in11[4];
    assign x11_5 = in11[5];
    assign x11_6 = in11[6];
    assign x11_7 = in11[7];
    assign x11_8 = in11[8];
    assign x11_9 = in11[9];
    assign x11_10 = in11[10];
    assign x11_11 = in11[11];
    assign x11_12 = in11[12];
    assign x11_13 = in11[13];
    assign x11_14 = in11[14];
    assign x11_15 = in11[15];
    assign x11_16 = in11[16];
    assign x11_17 = in11[17];
    assign x11_18 = in11[18];
    assign x11_19 = in11[19];
    assign x11_20 = in11[20];
    assign x11_21 = in11[21];
    assign x11_22 = in11[22];
    assign x11_23 = in11[23];
    assign x11_24 = in11[24];
    assign x11_25 = in11[25];
    assign x11_26 = in11[26];
    assign x11_27 = in11[27];
    assign x11_28 = in11[28];
    assign x11_29 = in11[29];
    assign x11_30 = in11[30];
    assign x11_31 = in11[31];
    assign x11_32 = in11[32];
    assign x11_33 = in11[33];
    assign x11_34 = in11[34];
    assign x11_35 = in11[35];
    assign x11_36 = in11[36];
    assign x11_37 = in11[37];
    assign x11_38 = in11[38];
    assign x11_39 = in11[39];
    assign x11_40 = in11[40];
    assign x11_41 = in11[41];
    assign x11_42 = in11[42];
    assign x11_43 = in11[43];
    assign x11_44 = in11[44];
    assign x11_45 = in11[45];
    assign x11_46 = in11[46];
    assign x11_47 = in11[47];
    assign x11_48 = in11[48];
    assign x11_49 = in11[49];
    assign x11_50 = in11[50];
    assign x11_51 = in11[51];
    assign x11_52 = in11[52];
    assign x11_53 = in11[53];
    assign x11_54 = in11[54];
    assign x11_55 = in11[55];
    assign x11_56 = in11[56];
    assign x11_57 = in11[57];
    assign x11_58 = in11[58];
    assign x11_59 = in11[59];
    assign x11_60 = in11[60];
    assign x11_61 = in11[61];
    assign x11_62 = in11[62];
    assign x11_63 = in11[63];
    assign x11_64 = in11[64];
    assign x11_65 = in11[65];
    assign x11_66 = in11[66];
    assign x11_67 = in11[67];
    assign x11_68 = in11[68];
    assign x11_69 = in11[69];
    wire x12_0;
    wire x12_1;
    wire x12_2;
    wire x12_3;
    wire x12_4;
    wire x12_5;
    wire x12_6;
    wire x12_7;
    wire x12_8;
    wire x12_9;
    wire x12_10;
    wire x12_11;
    wire x12_12;
    wire x12_13;
    wire x12_14;
    wire x12_15;
    wire x12_16;
    wire x12_17;
    wire x12_18;
    wire x12_19;
    wire x12_20;
    wire x12_21;
    wire x12_22;
    wire x12_23;
    wire x12_24;
    wire x12_25;
    wire x12_26;
    wire x12_27;
    wire x12_28;
    wire x12_29;
    wire x12_30;
    wire x12_31;
    wire x12_32;
    wire x12_33;
    wire x12_34;
    wire x12_35;
    wire x12_36;
    wire x12_37;
    wire x12_38;
    wire x12_39;
    wire x12_40;
    wire x12_41;
    wire x12_42;
    wire x12_43;
    wire x12_44;
    wire x12_45;
    wire x12_46;
    wire x12_47;
    wire x12_48;
    wire x12_49;
    wire x12_50;
    wire x12_51;
    wire x12_52;
    wire x12_53;
    wire x12_54;
    wire x12_55;
    wire x12_56;
    wire x12_57;
    wire x12_58;
    wire x12_59;
    wire x12_60;
    wire x12_61;
    wire x12_62;
    wire x12_63;
    wire x12_64;
    wire x12_65;
    wire x12_66;
    wire x12_67;
    wire x12_68;
    wire x12_69;
    assign x12_0 = in12[0];
    assign x12_1 = in12[1];
    assign x12_2 = in12[2];
    assign x12_3 = in12[3];
    assign x12_4 = in12[4];
    assign x12_5 = in12[5];
    assign x12_6 = in12[6];
    assign x12_7 = in12[7];
    assign x12_8 = in12[8];
    assign x12_9 = in12[9];
    assign x12_10 = in12[10];
    assign x12_11 = in12[11];
    assign x12_12 = in12[12];
    assign x12_13 = in12[13];
    assign x12_14 = in12[14];
    assign x12_15 = in12[15];
    assign x12_16 = in12[16];
    assign x12_17 = in12[17];
    assign x12_18 = in12[18];
    assign x12_19 = in12[19];
    assign x12_20 = in12[20];
    assign x12_21 = in12[21];
    assign x12_22 = in12[22];
    assign x12_23 = in12[23];
    assign x12_24 = in12[24];
    assign x12_25 = in12[25];
    assign x12_26 = in12[26];
    assign x12_27 = in12[27];
    assign x12_28 = in12[28];
    assign x12_29 = in12[29];
    assign x12_30 = in12[30];
    assign x12_31 = in12[31];
    assign x12_32 = in12[32];
    assign x12_33 = in12[33];
    assign x12_34 = in12[34];
    assign x12_35 = in12[35];
    assign x12_36 = in12[36];
    assign x12_37 = in12[37];
    assign x12_38 = in12[38];
    assign x12_39 = in12[39];
    assign x12_40 = in12[40];
    assign x12_41 = in12[41];
    assign x12_42 = in12[42];
    assign x12_43 = in12[43];
    assign x12_44 = in12[44];
    assign x12_45 = in12[45];
    assign x12_46 = in12[46];
    assign x12_47 = in12[47];
    assign x12_48 = in12[48];
    assign x12_49 = in12[49];
    assign x12_50 = in12[50];
    assign x12_51 = in12[51];
    assign x12_52 = in12[52];
    assign x12_53 = in12[53];
    assign x12_54 = in12[54];
    assign x12_55 = in12[55];
    assign x12_56 = in12[56];
    assign x12_57 = in12[57];
    assign x12_58 = in12[58];
    assign x12_59 = in12[59];
    assign x12_60 = in12[60];
    assign x12_61 = in12[61];
    assign x12_62 = in12[62];
    assign x12_63 = in12[63];
    assign x12_64 = in12[64];
    assign x12_65 = in12[65];
    assign x12_66 = in12[66];
    assign x12_67 = in12[67];
    assign x12_68 = in12[68];
    assign x12_69 = in12[69];
    wire x13_0;
    wire x13_1;
    wire x13_2;
    wire x13_3;
    wire x13_4;
    wire x13_5;
    wire x13_6;
    wire x13_7;
    wire x13_8;
    wire x13_9;
    wire x13_10;
    wire x13_11;
    wire x13_12;
    wire x13_13;
    wire x13_14;
    wire x13_15;
    wire x13_16;
    wire x13_17;
    wire x13_18;
    wire x13_19;
    wire x13_20;
    wire x13_21;
    wire x13_22;
    wire x13_23;
    wire x13_24;
    wire x13_25;
    wire x13_26;
    wire x13_27;
    wire x13_28;
    wire x13_29;
    wire x13_30;
    wire x13_31;
    wire x13_32;
    wire x13_33;
    wire x13_34;
    wire x13_35;
    wire x13_36;
    wire x13_37;
    wire x13_38;
    wire x13_39;
    wire x13_40;
    wire x13_41;
    wire x13_42;
    wire x13_43;
    wire x13_44;
    wire x13_45;
    wire x13_46;
    wire x13_47;
    wire x13_48;
    wire x13_49;
    wire x13_50;
    wire x13_51;
    wire x13_52;
    wire x13_53;
    wire x13_54;
    wire x13_55;
    wire x13_56;
    wire x13_57;
    wire x13_58;
    wire x13_59;
    wire x13_60;
    wire x13_61;
    wire x13_62;
    wire x13_63;
    wire x13_64;
    wire x13_65;
    wire x13_66;
    wire x13_67;
    wire x13_68;
    wire x13_69;
    assign x13_0 = in13[0];
    assign x13_1 = in13[1];
    assign x13_2 = in13[2];
    assign x13_3 = in13[3];
    assign x13_4 = in13[4];
    assign x13_5 = in13[5];
    assign x13_6 = in13[6];
    assign x13_7 = in13[7];
    assign x13_8 = in13[8];
    assign x13_9 = in13[9];
    assign x13_10 = in13[10];
    assign x13_11 = in13[11];
    assign x13_12 = in13[12];
    assign x13_13 = in13[13];
    assign x13_14 = in13[14];
    assign x13_15 = in13[15];
    assign x13_16 = in13[16];
    assign x13_17 = in13[17];
    assign x13_18 = in13[18];
    assign x13_19 = in13[19];
    assign x13_20 = in13[20];
    assign x13_21 = in13[21];
    assign x13_22 = in13[22];
    assign x13_23 = in13[23];
    assign x13_24 = in13[24];
    assign x13_25 = in13[25];
    assign x13_26 = in13[26];
    assign x13_27 = in13[27];
    assign x13_28 = in13[28];
    assign x13_29 = in13[29];
    assign x13_30 = in13[30];
    assign x13_31 = in13[31];
    assign x13_32 = in13[32];
    assign x13_33 = in13[33];
    assign x13_34 = in13[34];
    assign x13_35 = in13[35];
    assign x13_36 = in13[36];
    assign x13_37 = in13[37];
    assign x13_38 = in13[38];
    assign x13_39 = in13[39];
    assign x13_40 = in13[40];
    assign x13_41 = in13[41];
    assign x13_42 = in13[42];
    assign x13_43 = in13[43];
    assign x13_44 = in13[44];
    assign x13_45 = in13[45];
    assign x13_46 = in13[46];
    assign x13_47 = in13[47];
    assign x13_48 = in13[48];
    assign x13_49 = in13[49];
    assign x13_50 = in13[50];
    assign x13_51 = in13[51];
    assign x13_52 = in13[52];
    assign x13_53 = in13[53];
    assign x13_54 = in13[54];
    assign x13_55 = in13[55];
    assign x13_56 = in13[56];
    assign x13_57 = in13[57];
    assign x13_58 = in13[58];
    assign x13_59 = in13[59];
    assign x13_60 = in13[60];
    assign x13_61 = in13[61];
    assign x13_62 = in13[62];
    assign x13_63 = in13[63];
    assign x13_64 = in13[64];
    assign x13_65 = in13[65];
    assign x13_66 = in13[66];
    assign x13_67 = in13[67];
    assign x13_68 = in13[68];
    assign x13_69 = in13[69];
    wire x14_0;
    wire x14_1;
    wire x14_2;
    wire x14_3;
    wire x14_4;
    wire x14_5;
    wire x14_6;
    wire x14_7;
    wire x14_8;
    wire x14_9;
    wire x14_10;
    wire x14_11;
    wire x14_12;
    wire x14_13;
    wire x14_14;
    wire x14_15;
    wire x14_16;
    wire x14_17;
    wire x14_18;
    wire x14_19;
    wire x14_20;
    wire x14_21;
    wire x14_22;
    wire x14_23;
    wire x14_24;
    wire x14_25;
    wire x14_26;
    wire x14_27;
    wire x14_28;
    wire x14_29;
    wire x14_30;
    wire x14_31;
    wire x14_32;
    wire x14_33;
    wire x14_34;
    wire x14_35;
    wire x14_36;
    wire x14_37;
    wire x14_38;
    wire x14_39;
    wire x14_40;
    wire x14_41;
    wire x14_42;
    wire x14_43;
    wire x14_44;
    wire x14_45;
    wire x14_46;
    wire x14_47;
    wire x14_48;
    wire x14_49;
    wire x14_50;
    wire x14_51;
    wire x14_52;
    wire x14_53;
    wire x14_54;
    wire x14_55;
    wire x14_56;
    wire x14_57;
    wire x14_58;
    wire x14_59;
    wire x14_60;
    wire x14_61;
    wire x14_62;
    wire x14_63;
    wire x14_64;
    wire x14_65;
    wire x14_66;
    wire x14_67;
    wire x14_68;
    wire x14_69;
    assign x14_0 = in14[0];
    assign x14_1 = in14[1];
    assign x14_2 = in14[2];
    assign x14_3 = in14[3];
    assign x14_4 = in14[4];
    assign x14_5 = in14[5];
    assign x14_6 = in14[6];
    assign x14_7 = in14[7];
    assign x14_8 = in14[8];
    assign x14_9 = in14[9];
    assign x14_10 = in14[10];
    assign x14_11 = in14[11];
    assign x14_12 = in14[12];
    assign x14_13 = in14[13];
    assign x14_14 = in14[14];
    assign x14_15 = in14[15];
    assign x14_16 = in14[16];
    assign x14_17 = in14[17];
    assign x14_18 = in14[18];
    assign x14_19 = in14[19];
    assign x14_20 = in14[20];
    assign x14_21 = in14[21];
    assign x14_22 = in14[22];
    assign x14_23 = in14[23];
    assign x14_24 = in14[24];
    assign x14_25 = in14[25];
    assign x14_26 = in14[26];
    assign x14_27 = in14[27];
    assign x14_28 = in14[28];
    assign x14_29 = in14[29];
    assign x14_30 = in14[30];
    assign x14_31 = in14[31];
    assign x14_32 = in14[32];
    assign x14_33 = in14[33];
    assign x14_34 = in14[34];
    assign x14_35 = in14[35];
    assign x14_36 = in14[36];
    assign x14_37 = in14[37];
    assign x14_38 = in14[38];
    assign x14_39 = in14[39];
    assign x14_40 = in14[40];
    assign x14_41 = in14[41];
    assign x14_42 = in14[42];
    assign x14_43 = in14[43];
    assign x14_44 = in14[44];
    assign x14_45 = in14[45];
    assign x14_46 = in14[46];
    assign x14_47 = in14[47];
    assign x14_48 = in14[48];
    assign x14_49 = in14[49];
    assign x14_50 = in14[50];
    assign x14_51 = in14[51];
    assign x14_52 = in14[52];
    assign x14_53 = in14[53];
    assign x14_54 = in14[54];
    assign x14_55 = in14[55];
    assign x14_56 = in14[56];
    assign x14_57 = in14[57];
    assign x14_58 = in14[58];
    assign x14_59 = in14[59];
    assign x14_60 = in14[60];
    assign x14_61 = in14[61];
    assign x14_62 = in14[62];
    assign x14_63 = in14[63];
    assign x14_64 = in14[64];
    assign x14_65 = in14[65];
    assign x14_66 = in14[66];
    assign x14_67 = in14[67];
    assign x14_68 = in14[68];
    assign x14_69 = in14[69];
    wire x15_0;
    wire x15_1;
    wire x15_2;
    wire x15_3;
    wire x15_4;
    wire x15_5;
    wire x15_6;
    wire x15_7;
    wire x15_8;
    wire x15_9;
    wire x15_10;
    wire x15_11;
    wire x15_12;
    wire x15_13;
    wire x15_14;
    wire x15_15;
    wire x15_16;
    wire x15_17;
    wire x15_18;
    wire x15_19;
    wire x15_20;
    wire x15_21;
    wire x15_22;
    wire x15_23;
    wire x15_24;
    wire x15_25;
    wire x15_26;
    wire x15_27;
    wire x15_28;
    wire x15_29;
    wire x15_30;
    wire x15_31;
    wire x15_32;
    wire x15_33;
    wire x15_34;
    wire x15_35;
    wire x15_36;
    wire x15_37;
    wire x15_38;
    wire x15_39;
    wire x15_40;
    wire x15_41;
    wire x15_42;
    wire x15_43;
    wire x15_44;
    wire x15_45;
    wire x15_46;
    wire x15_47;
    wire x15_48;
    wire x15_49;
    wire x15_50;
    wire x15_51;
    wire x15_52;
    wire x15_53;
    wire x15_54;
    wire x15_55;
    wire x15_56;
    wire x15_57;
    wire x15_58;
    wire x15_59;
    wire x15_60;
    wire x15_61;
    wire x15_62;
    wire x15_63;
    wire x15_64;
    wire x15_65;
    wire x15_66;
    wire x15_67;
    wire x15_68;
    wire x15_69;
    assign x15_0 = in15[0];
    assign x15_1 = in15[1];
    assign x15_2 = in15[2];
    assign x15_3 = in15[3];
    assign x15_4 = in15[4];
    assign x15_5 = in15[5];
    assign x15_6 = in15[6];
    assign x15_7 = in15[7];
    assign x15_8 = in15[8];
    assign x15_9 = in15[9];
    assign x15_10 = in15[10];
    assign x15_11 = in15[11];
    assign x15_12 = in15[12];
    assign x15_13 = in15[13];
    assign x15_14 = in15[14];
    assign x15_15 = in15[15];
    assign x15_16 = in15[16];
    assign x15_17 = in15[17];
    assign x15_18 = in15[18];
    assign x15_19 = in15[19];
    assign x15_20 = in15[20];
    assign x15_21 = in15[21];
    assign x15_22 = in15[22];
    assign x15_23 = in15[23];
    assign x15_24 = in15[24];
    assign x15_25 = in15[25];
    assign x15_26 = in15[26];
    assign x15_27 = in15[27];
    assign x15_28 = in15[28];
    assign x15_29 = in15[29];
    assign x15_30 = in15[30];
    assign x15_31 = in15[31];
    assign x15_32 = in15[32];
    assign x15_33 = in15[33];
    assign x15_34 = in15[34];
    assign x15_35 = in15[35];
    assign x15_36 = in15[36];
    assign x15_37 = in15[37];
    assign x15_38 = in15[38];
    assign x15_39 = in15[39];
    assign x15_40 = in15[40];
    assign x15_41 = in15[41];
    assign x15_42 = in15[42];
    assign x15_43 = in15[43];
    assign x15_44 = in15[44];
    assign x15_45 = in15[45];
    assign x15_46 = in15[46];
    assign x15_47 = in15[47];
    assign x15_48 = in15[48];
    assign x15_49 = in15[49];
    assign x15_50 = in15[50];
    assign x15_51 = in15[51];
    assign x15_52 = in15[52];
    assign x15_53 = in15[53];
    assign x15_54 = in15[54];
    assign x15_55 = in15[55];
    assign x15_56 = in15[56];
    assign x15_57 = in15[57];
    assign x15_58 = in15[58];
    assign x15_59 = in15[59];
    assign x15_60 = in15[60];
    assign x15_61 = in15[61];
    assign x15_62 = in15[62];
    assign x15_63 = in15[63];
    assign x15_64 = in15[64];
    assign x15_65 = in15[65];
    assign x15_66 = in15[66];
    assign x15_67 = in15[67];
    assign x15_68 = in15[68];
    assign x15_69 = in15[69];
    wire w1;
    wire w2;
    wire w3;
    wire w4;
    wire w5;
    wire w6;
    wire w7;
    wire w8;
    wire w9;
    wire w10;
    wire w11;
    wire w12;
    wire w13;
    wire w14;
    wire w15;
    wire w16;
    wire w17;
    wire w18;
    wire w19;
    wire w20;
    wire w21;
    wire w22;
    wire w23;
    wire w24;
    wire w25;
    wire w26;
    wire w27;
    wire w28;
    wire w29;
    wire w30;
    wire w31;
    wire w32;
    wire w33;
    wire w34;
    wire w35;
    wire w36;
    wire w37;
    wire w38;
    wire w39;
    wire w40;
    wire w41;
    wire w42;
    wire w43;
    wire w44;
    wire w45;
    wire w46;
    wire w47;
    wire w48;
    wire w49;
    wire w50;
    wire w51;
    wire w52;
    wire w53;
    wire w54;
    wire w55;
    wire w56;
    wire w57;
    wire w58;
    wire w59;
    wire w60;
    wire w61;
    wire w62;
    wire w63;
    wire w64;
    wire w65;
    wire w66;
    wire w67;
    wire w68;
    wire w69;
    assign out0[0] = w1;
    assign out0[1] = w2;
    assign out0[2] = w3;
    assign out0[3] = w4;
    assign out0[4] = w5;
    assign out0[5] = w6;
    assign out0[6] = w7;
    assign out0[7] = w8;
    assign out0[8] = w9;
    assign out0[9] = w10;
    assign out0[10] = w11;
    assign out0[11] = w12;
    assign out0[12] = w13;
    assign out0[13] = w14;
    assign out0[14] = w15;
    assign out0[15] = w16;
    assign out0[16] = w17;
    assign out0[17] = w18;
    assign out0[18] = w19;
    assign out0[19] = w20;
    assign out0[20] = w21;
    assign out0[21] = w22;
    assign out0[22] = w23;
    assign out0[23] = w24;
    assign out0[24] = w25;
    assign out0[25] = w26;
    assign out0[26] = w27;
    assign out0[27] = w28;
    assign out0[28] = w29;
    assign out0[29] = w30;
    assign out0[30] = w31;
    assign out0[31] = w32;
    assign out0[32] = w33;
    assign out0[33] = w34;
    assign out0[34] = w35;
    assign out0[35] = w36;
    assign out0[36] = w37;
    assign out0[37] = w38;
    assign out0[38] = w39;
    assign out0[39] = w40;
    assign out0[40] = w41;
    assign out0[41] = w42;
    assign out0[42] = w43;
    assign out0[43] = w44;
    assign out0[44] = w45;
    assign out0[45] = w46;
    assign out0[46] = w47;
    assign out0[47] = w48;
    assign out0[48] = w49;
    assign out0[49] = w50;
    assign out0[50] = w51;
    assign out0[51] = w52;
    assign out0[52] = w53;
    assign out0[53] = w54;
    assign out0[54] = w55;
    assign out0[55] = w56;
    assign out0[56] = w57;
    assign out0[57] = w58;
    assign out0[58] = w59;
    assign out0[59] = w60;
    assign out0[60] = w61;
    assign out0[61] = w62;
    assign out0[62] = w63;
    assign out0[63] = w64;
    assign out0[64] = w65;
    assign out0[65] = w66;
    assign out0[66] = w67;
    assign out0[67] = w68;
    assign out0[68] = w69;
    wire w70;
    wire w71;
    wire w72;
    wire w73;
    wire w74;
    wire w75;
    wire w76;
    wire w77;
    wire w78;
    wire w79;
    wire w80;
    wire w81;
    wire w82;
    wire w83;
    wire w84;
    wire w85;
    wire w86;
    wire w87;
    wire w88;
    wire w89;
    wire w90;
    wire w91;
    wire w92;
    wire w93;
    wire w94;
    wire w95;
    wire w96;
    wire w97;
    wire w98;
    wire w99;
    wire w100;
    wire w101;
    wire w102;
    wire w103;
    wire w104;
    wire w105;
    wire w106;
    wire w107;
    wire w108;
    wire w109;
    wire w110;
    wire w111;
    wire w112;
    wire w113;
    wire w114;
    wire w115;
    wire w116;
    wire w117;
    wire w118;
    wire w119;
    wire w120;
    wire w121;
    wire w122;
    wire w123;
    wire w124;
    wire w125;
    wire w126;
    wire w127;
    wire w128;
    wire w129;
    wire w130;
    wire w131;
    wire w132;
    wire w133;
    wire w134;
    wire w135;
    wire w136;
    wire w137;
    wire w138;
    assign out1[0] = w70;
    assign out1[1] = w71;
    assign out1[2] = w72;
    assign out1[3] = w73;
    assign out1[4] = w74;
    assign out1[5] = w75;
    assign out1[6] = w76;
    assign out1[7] = w77;
    assign out1[8] = w78;
    assign out1[9] = w79;
    assign out1[10] = w80;
    assign out1[11] = w81;
    assign out1[12] = w82;
    assign out1[13] = w83;
    assign out1[14] = w84;
    assign out1[15] = w85;
    assign out1[16] = w86;
    assign out1[17] = w87;
    assign out1[18] = w88;
    assign out1[19] = w89;
    assign out1[20] = w90;
    assign out1[21] = w91;
    assign out1[22] = w92;
    assign out1[23] = w93;
    assign out1[24] = w94;
    assign out1[25] = w95;
    assign out1[26] = w96;
    assign out1[27] = w97;
    assign out1[28] = w98;
    assign out1[29] = w99;
    assign out1[30] = w100;
    assign out1[31] = w101;
    assign out1[32] = w102;
    assign out1[33] = w103;
    assign out1[34] = w104;
    assign out1[35] = w105;
    assign out1[36] = w106;
    assign out1[37] = w107;
    assign out1[38] = w108;
    assign out1[39] = w109;
    assign out1[40] = w110;
    assign out1[41] = w111;
    assign out1[42] = w112;
    assign out1[43] = w113;
    assign out1[44] = w114;
    assign out1[45] = w115;
    assign out1[46] = w116;
    assign out1[47] = w117;
    assign out1[48] = w118;
    assign out1[49] = w119;
    assign out1[50] = w120;
    assign out1[51] = w121;
    assign out1[52] = w122;
    assign out1[53] = w123;
    assign out1[54] = w124;
    assign out1[55] = w125;
    assign out1[56] = w126;
    assign out1[57] = w127;
    assign out1[58] = w128;
    assign out1[59] = w129;
    assign out1[60] = w130;
    assign out1[61] = w131;
    assign out1[62] = w132;
    assign out1[63] = w133;
    assign out1[64] = w134;
    assign out1[65] = w135;
    assign out1[66] = w136;
    assign out1[67] = w137;
    assign out1[68] = w138;
    wire w139;
    wire w140;
    wire w141;
    wire w142;
    wire w143;
    wire w144;
    wire w145;
    wire w146;
    wire w147;
    wire w148;
    wire w149;
    wire w150;
    wire w151;
    wire w152;
    wire w153;
    wire w154;
    wire w155;
    wire w156;
    wire w157;
    wire w158;
    wire w159;
    wire w160;
    wire w161;
    wire w162;
    wire w163;
    wire w164;
    wire w165;
    wire w166;
    wire w167;
    wire w168;
    wire w169;
    wire w170;
    wire w171;
    wire w172;
    wire w173;
    wire w174;
    wire w175;
    wire w176;
    wire w177;
    wire w178;
    wire w179;
    wire w180;
    wire w181;
    wire w182;
    wire w183;
    wire w184;
    wire w185;
    wire w186;
    wire w187;
    wire w188;
    wire w189;
    wire w190;
    wire w191;
    wire w192;
    wire w193;
    wire w194;
    wire w195;
    wire w196;
    wire w197;
    wire w198;
    wire w199;
    wire w200;
    wire w201;
    wire w202;
    wire w203;
    wire w204;
    wire w205;
    wire w206;
    wire w207;
    assign out2[0] = w139;
    assign out2[1] = w140;
    assign out2[2] = w141;
    assign out2[3] = w142;
    assign out2[4] = w143;
    assign out2[5] = w144;
    assign out2[6] = w145;
    assign out2[7] = w146;
    assign out2[8] = w147;
    assign out2[9] = w148;
    assign out2[10] = w149;
    assign out2[11] = w150;
    assign out2[12] = w151;
    assign out2[13] = w152;
    assign out2[14] = w153;
    assign out2[15] = w154;
    assign out2[16] = w155;
    assign out2[17] = w156;
    assign out2[18] = w157;
    assign out2[19] = w158;
    assign out2[20] = w159;
    assign out2[21] = w160;
    assign out2[22] = w161;
    assign out2[23] = w162;
    assign out2[24] = w163;
    assign out2[25] = w164;
    assign out2[26] = w165;
    assign out2[27] = w166;
    assign out2[28] = w167;
    assign out2[29] = w168;
    assign out2[30] = w169;
    assign out2[31] = w170;
    assign out2[32] = w171;
    assign out2[33] = w172;
    assign out2[34] = w173;
    assign out2[35] = w174;
    assign out2[36] = w175;
    assign out2[37] = w176;
    assign out2[38] = w177;
    assign out2[39] = w178;
    assign out2[40] = w179;
    assign out2[41] = w180;
    assign out2[42] = w181;
    assign out2[43] = w182;
    assign out2[44] = w183;
    assign out2[45] = w184;
    assign out2[46] = w185;
    assign out2[47] = w186;
    assign out2[48] = w187;
    assign out2[49] = w188;
    assign out2[50] = w189;
    assign out2[51] = w190;
    assign out2[52] = w191;
    assign out2[53] = w192;
    assign out2[54] = w193;
    assign out2[55] = w194;
    assign out2[56] = w195;
    assign out2[57] = w196;
    assign out2[58] = w197;
    assign out2[59] = w198;
    assign out2[60] = w199;
    assign out2[61] = w200;
    assign out2[62] = w201;
    assign out2[63] = w202;
    assign out2[64] = w203;
    assign out2[65] = w204;
    assign out2[66] = w205;
    assign out2[67] = w206;
    assign out2[68] = w207;
    wire w208;
    wire w209;
    wire w210;
    wire w211;
    wire w212;
    wire w213;
    wire w214;
    wire w215;
    wire w216;
    wire w217;
    wire w218;
    wire w219;
    wire w220;
    wire w221;
    wire w222;
    wire w223;
    wire w224;
    wire w225;
    wire w226;
    wire w227;
    wire w228;
    wire w229;
    wire w230;
    wire w231;
    wire w232;
    wire w233;
    wire w234;
    wire w235;
    wire w236;
    wire w237;
    wire w238;
    wire w239;
    wire w240;
    wire w241;
    wire w242;
    wire w243;
    wire w244;
    wire w245;
    wire w246;
    wire w247;
    wire w248;
    wire w249;
    wire w250;
    wire w251;
    wire w252;
    wire w253;
    wire w254;
    wire w255;
    wire w256;
    wire w257;
    wire w258;
    wire w259;
    wire w260;
    wire w261;
    wire w262;
    wire w263;
    wire w264;
    wire w265;
    wire w266;
    wire w267;
    wire w268;
    wire w269;
    wire w270;
    wire w271;
    wire w272;
    wire w273;
    wire w274;
    wire w275;
    wire w276;
    assign out3[0] = w208;
    assign out3[1] = w209;
    assign out3[2] = w210;
    assign out3[3] = w211;
    assign out3[4] = w212;
    assign out3[5] = w213;
    assign out3[6] = w214;
    assign out3[7] = w215;
    assign out3[8] = w216;
    assign out3[9] = w217;
    assign out3[10] = w218;
    assign out3[11] = w219;
    assign out3[12] = w220;
    assign out3[13] = w221;
    assign out3[14] = w222;
    assign out3[15] = w223;
    assign out3[16] = w224;
    assign out3[17] = w225;
    assign out3[18] = w226;
    assign out3[19] = w227;
    assign out3[20] = w228;
    assign out3[21] = w229;
    assign out3[22] = w230;
    assign out3[23] = w231;
    assign out3[24] = w232;
    assign out3[25] = w233;
    assign out3[26] = w234;
    assign out3[27] = w235;
    assign out3[28] = w236;
    assign out3[29] = w237;
    assign out3[30] = w238;
    assign out3[31] = w239;
    assign out3[32] = w240;
    assign out3[33] = w241;
    assign out3[34] = w242;
    assign out3[35] = w243;
    assign out3[36] = w244;
    assign out3[37] = w245;
    assign out3[38] = w246;
    assign out3[39] = w247;
    assign out3[40] = w248;
    assign out3[41] = w249;
    assign out3[42] = w250;
    assign out3[43] = w251;
    assign out3[44] = w252;
    assign out3[45] = w253;
    assign out3[46] = w254;
    assign out3[47] = w255;
    assign out3[48] = w256;
    assign out3[49] = w257;
    assign out3[50] = w258;
    assign out3[51] = w259;
    assign out3[52] = w260;
    assign out3[53] = w261;
    assign out3[54] = w262;
    assign out3[55] = w263;
    assign out3[56] = w264;
    assign out3[57] = w265;
    assign out3[58] = w266;
    assign out3[59] = w267;
    assign out3[60] = w268;
    assign out3[61] = w269;
    assign out3[62] = w270;
    assign out3[63] = w271;
    assign out3[64] = w272;
    assign out3[65] = w273;
    assign out3[66] = w274;
    assign out3[67] = w275;
    assign out3[68] = w276;
    wire w277;
    wire w278;
    wire w279;
    wire w280;
    wire w281;
    wire w282;
    wire w283;
    wire w284;
    wire w285;
    wire w286;
    wire w287;
    wire w288;
    wire w289;
    wire w290;
    wire w291;
    wire w292;
    wire w293;
    wire w294;
    wire w295;
    wire w296;
    wire w297;
    wire w298;
    wire w299;
    wire w300;
    wire w301;
    wire w302;
    wire w303;
    wire w304;
    wire w305;
    wire w306;
    wire w307;
    wire w308;
    wire w309;
    wire w310;
    wire w311;
    wire w312;
    wire w313;
    wire w314;
    wire w315;
    wire w316;
    wire w317;
    wire w318;
    wire w319;
    wire w320;
    wire w321;
    wire w322;
    wire w323;
    wire w324;
    wire w325;
    wire w326;
    wire w327;
    wire w328;
    wire w329;
    wire w330;
    wire w331;
    wire w332;
    wire w333;
    wire w334;
    wire w335;
    wire w336;
    wire w337;
    wire w338;
    wire w339;
    wire w340;
    wire w341;
    wire w342;
    wire w343;
    wire w344;
    wire w345;
    assign out4[0] = w277;
    assign out4[1] = w278;
    assign out4[2] = w279;
    assign out4[3] = w280;
    assign out4[4] = w281;
    assign out4[5] = w282;
    assign out4[6] = w283;
    assign out4[7] = w284;
    assign out4[8] = w285;
    assign out4[9] = w286;
    assign out4[10] = w287;
    assign out4[11] = w288;
    assign out4[12] = w289;
    assign out4[13] = w290;
    assign out4[14] = w291;
    assign out4[15] = w292;
    assign out4[16] = w293;
    assign out4[17] = w294;
    assign out4[18] = w295;
    assign out4[19] = w296;
    assign out4[20] = w297;
    assign out4[21] = w298;
    assign out4[22] = w299;
    assign out4[23] = w300;
    assign out4[24] = w301;
    assign out4[25] = w302;
    assign out4[26] = w303;
    assign out4[27] = w304;
    assign out4[28] = w305;
    assign out4[29] = w306;
    assign out4[30] = w307;
    assign out4[31] = w308;
    assign out4[32] = w309;
    assign out4[33] = w310;
    assign out4[34] = w311;
    assign out4[35] = w312;
    assign out4[36] = w313;
    assign out4[37] = w314;
    assign out4[38] = w315;
    assign out4[39] = w316;
    assign out4[40] = w317;
    assign out4[41] = w318;
    assign out4[42] = w319;
    assign out4[43] = w320;
    assign out4[44] = w321;
    assign out4[45] = w322;
    assign out4[46] = w323;
    assign out4[47] = w324;
    assign out4[48] = w325;
    assign out4[49] = w326;
    assign out4[50] = w327;
    assign out4[51] = w328;
    assign out4[52] = w329;
    assign out4[53] = w330;
    assign out4[54] = w331;
    assign out4[55] = w332;
    assign out4[56] = w333;
    assign out4[57] = w334;
    assign out4[58] = w335;
    assign out4[59] = w336;
    assign out4[60] = w337;
    assign out4[61] = w338;
    assign out4[62] = w339;
    assign out4[63] = w340;
    assign out4[64] = w341;
    assign out4[65] = w342;
    assign out4[66] = w343;
    assign out4[67] = w344;
    assign out4[68] = w345;
    wire w346;
    wire w347;
    wire w348;
    wire w349;
    wire w350;
    wire w351;
    wire w352;
    wire w353;
    wire w354;
    wire w355;
    wire w356;
    wire w357;
    wire w358;
    wire w359;
    wire w360;
    wire w361;
    wire w362;
    wire w363;
    wire w364;
    wire w365;
    wire w366;
    wire w367;
    wire w368;
    wire w369;
    wire w370;
    wire w371;
    wire w372;
    wire w373;
    wire w374;
    wire w375;
    wire w376;
    wire w377;
    wire w378;
    wire w379;
    wire w380;
    wire w381;
    wire w382;
    wire w383;
    wire w384;
    wire w385;
    wire w386;
    wire w387;
    wire w388;
    wire w389;
    wire w390;
    wire w391;
    wire w392;
    wire w393;
    wire w394;
    wire w395;
    wire w396;
    wire w397;
    wire w398;
    wire w399;
    wire w400;
    wire w401;
    wire w402;
    wire w403;
    wire w404;
    wire w405;
    wire w406;
    wire w407;
    wire w408;
    wire w409;
    wire w410;
    wire w411;
    wire w412;
    wire w413;
    wire w414;
    assign out5[0] = w346;
    assign out5[1] = w347;
    assign out5[2] = w348;
    assign out5[3] = w349;
    assign out5[4] = w350;
    assign out5[5] = w351;
    assign out5[6] = w352;
    assign out5[7] = w353;
    assign out5[8] = w354;
    assign out5[9] = w355;
    assign out5[10] = w356;
    assign out5[11] = w357;
    assign out5[12] = w358;
    assign out5[13] = w359;
    assign out5[14] = w360;
    assign out5[15] = w361;
    assign out5[16] = w362;
    assign out5[17] = w363;
    assign out5[18] = w364;
    assign out5[19] = w365;
    assign out5[20] = w366;
    assign out5[21] = w367;
    assign out5[22] = w368;
    assign out5[23] = w369;
    assign out5[24] = w370;
    assign out5[25] = w371;
    assign out5[26] = w372;
    assign out5[27] = w373;
    assign out5[28] = w374;
    assign out5[29] = w375;
    assign out5[30] = w376;
    assign out5[31] = w377;
    assign out5[32] = w378;
    assign out5[33] = w379;
    assign out5[34] = w380;
    assign out5[35] = w381;
    assign out5[36] = w382;
    assign out5[37] = w383;
    assign out5[38] = w384;
    assign out5[39] = w385;
    assign out5[40] = w386;
    assign out5[41] = w387;
    assign out5[42] = w388;
    assign out5[43] = w389;
    assign out5[44] = w390;
    assign out5[45] = w391;
    assign out5[46] = w392;
    assign out5[47] = w393;
    assign out5[48] = w394;
    assign out5[49] = w395;
    assign out5[50] = w396;
    assign out5[51] = w397;
    assign out5[52] = w398;
    assign out5[53] = w399;
    assign out5[54] = w400;
    assign out5[55] = w401;
    assign out5[56] = w402;
    assign out5[57] = w403;
    assign out5[58] = w404;
    assign out5[59] = w405;
    assign out5[60] = w406;
    assign out5[61] = w407;
    assign out5[62] = w408;
    assign out5[63] = w409;
    assign out5[64] = w410;
    assign out5[65] = w411;
    assign out5[66] = w412;
    assign out5[67] = w413;
    assign out5[68] = w414;
    wire w415;
    wire w416;
    wire w417;
    wire w418;
    wire w419;
    wire w420;
    wire w421;
    wire w422;
    wire w423;
    wire w424;
    wire w425;
    wire w426;
    wire w427;
    wire w428;
    wire w429;
    wire w430;
    wire w431;
    wire w432;
    wire w433;
    wire w434;
    wire w435;
    wire w436;
    wire w437;
    wire w438;
    wire w439;
    wire w440;
    wire w441;
    wire w442;
    wire w443;
    wire w444;
    wire w445;
    wire w446;
    wire w447;
    wire w448;
    wire w449;
    wire w450;
    wire w451;
    wire w452;
    wire w453;
    wire w454;
    wire w455;
    wire w456;
    wire w457;
    wire w458;
    wire w459;
    wire w460;
    wire w461;
    wire w462;
    wire w463;
    wire w464;
    wire w465;
    wire w466;
    wire w467;
    wire w468;
    wire w469;
    wire w470;
    wire w471;
    wire w472;
    wire w473;
    wire w474;
    wire w475;
    wire w476;
    wire w477;
    wire w478;
    wire w479;
    wire w480;
    wire w481;
    wire w482;
    wire w483;
    assign out6[0] = w415;
    assign out6[1] = w416;
    assign out6[2] = w417;
    assign out6[3] = w418;
    assign out6[4] = w419;
    assign out6[5] = w420;
    assign out6[6] = w421;
    assign out6[7] = w422;
    assign out6[8] = w423;
    assign out6[9] = w424;
    assign out6[10] = w425;
    assign out6[11] = w426;
    assign out6[12] = w427;
    assign out6[13] = w428;
    assign out6[14] = w429;
    assign out6[15] = w430;
    assign out6[16] = w431;
    assign out6[17] = w432;
    assign out6[18] = w433;
    assign out6[19] = w434;
    assign out6[20] = w435;
    assign out6[21] = w436;
    assign out6[22] = w437;
    assign out6[23] = w438;
    assign out6[24] = w439;
    assign out6[25] = w440;
    assign out6[26] = w441;
    assign out6[27] = w442;
    assign out6[28] = w443;
    assign out6[29] = w444;
    assign out6[30] = w445;
    assign out6[31] = w446;
    assign out6[32] = w447;
    assign out6[33] = w448;
    assign out6[34] = w449;
    assign out6[35] = w450;
    assign out6[36] = w451;
    assign out6[37] = w452;
    assign out6[38] = w453;
    assign out6[39] = w454;
    assign out6[40] = w455;
    assign out6[41] = w456;
    assign out6[42] = w457;
    assign out6[43] = w458;
    assign out6[44] = w459;
    assign out6[45] = w460;
    assign out6[46] = w461;
    assign out6[47] = w462;
    assign out6[48] = w463;
    assign out6[49] = w464;
    assign out6[50] = w465;
    assign out6[51] = w466;
    assign out6[52] = w467;
    assign out6[53] = w468;
    assign out6[54] = w469;
    assign out6[55] = w470;
    assign out6[56] = w471;
    assign out6[57] = w472;
    assign out6[58] = w473;
    assign out6[59] = w474;
    assign out6[60] = w475;
    assign out6[61] = w476;
    assign out6[62] = w477;
    assign out6[63] = w478;
    assign out6[64] = w479;
    assign out6[65] = w480;
    assign out6[66] = w481;
    assign out6[67] = w482;
    assign out6[68] = w483;
    wire w484;
    wire w485;
    wire w486;
    wire w487;
    wire w488;
    wire w489;
    wire w490;
    wire w491;
    wire w492;
    wire w493;
    wire w494;
    wire w495;
    wire w496;
    wire w497;
    wire w498;
    wire w499;
    wire w500;
    wire w501;
    wire w502;
    wire w503;
    wire w504;
    wire w505;
    wire w506;
    wire w507;
    wire w508;
    wire w509;
    wire w510;
    wire w511;
    wire w512;
    wire w513;
    wire w514;
    wire w515;
    wire w516;
    wire w517;
    wire w518;
    wire w519;
    wire w520;
    wire w521;
    wire w522;
    wire w523;
    wire w524;
    wire w525;
    wire w526;
    wire w527;
    wire w528;
    wire w529;
    wire w530;
    wire w531;
    wire w532;
    wire w533;
    wire w534;
    wire w535;
    wire w536;
    wire w537;
    wire w538;
    wire w539;
    wire w540;
    wire w541;
    wire w542;
    wire w543;
    wire w544;
    wire w545;
    wire w546;
    wire w547;
    wire w548;
    wire w549;
    wire w550;
    wire w551;
    wire w552;
    assign out7[0] = w484;
    assign out7[1] = w485;
    assign out7[2] = w486;
    assign out7[3] = w487;
    assign out7[4] = w488;
    assign out7[5] = w489;
    assign out7[6] = w490;
    assign out7[7] = w491;
    assign out7[8] = w492;
    assign out7[9] = w493;
    assign out7[10] = w494;
    assign out7[11] = w495;
    assign out7[12] = w496;
    assign out7[13] = w497;
    assign out7[14] = w498;
    assign out7[15] = w499;
    assign out7[16] = w500;
    assign out7[17] = w501;
    assign out7[18] = w502;
    assign out7[19] = w503;
    assign out7[20] = w504;
    assign out7[21] = w505;
    assign out7[22] = w506;
    assign out7[23] = w507;
    assign out7[24] = w508;
    assign out7[25] = w509;
    assign out7[26] = w510;
    assign out7[27] = w511;
    assign out7[28] = w512;
    assign out7[29] = w513;
    assign out7[30] = w514;
    assign out7[31] = w515;
    assign out7[32] = w516;
    assign out7[33] = w517;
    assign out7[34] = w518;
    assign out7[35] = w519;
    assign out7[36] = w520;
    assign out7[37] = w521;
    assign out7[38] = w522;
    assign out7[39] = w523;
    assign out7[40] = w524;
    assign out7[41] = w525;
    assign out7[42] = w526;
    assign out7[43] = w527;
    assign out7[44] = w528;
    assign out7[45] = w529;
    assign out7[46] = w530;
    assign out7[47] = w531;
    assign out7[48] = w532;
    assign out7[49] = w533;
    assign out7[50] = w534;
    assign out7[51] = w535;
    assign out7[52] = w536;
    assign out7[53] = w537;
    assign out7[54] = w538;
    assign out7[55] = w539;
    assign out7[56] = w540;
    assign out7[57] = w541;
    assign out7[58] = w542;
    assign out7[59] = w543;
    assign out7[60] = w544;
    assign out7[61] = w545;
    assign out7[62] = w546;
    assign out7[63] = w547;
    assign out7[64] = w548;
    assign out7[65] = w549;
    assign out7[66] = w550;
    assign out7[67] = w551;
    assign out7[68] = w552;
    wire w553;
    wire w554;
    wire w555;
    wire w556;
    wire w557;
    wire w558;
    wire w559;
    wire w560;
    wire w561;
    wire w562;
    wire w563;
    wire w564;
    wire w565;
    wire w566;
    wire w567;
    wire w568;
    wire w569;
    wire w570;
    wire w571;
    wire w572;
    wire w573;
    wire w574;
    wire w575;
    wire w576;
    wire w577;
    wire w578;
    wire w579;
    wire w580;
    wire w581;
    wire w582;
    wire w583;
    wire w584;
    wire w585;
    wire w586;
    wire w587;
    wire w588;
    wire w589;
    wire w590;
    wire w591;
    wire w592;
    wire w593;
    wire w594;
    wire w595;
    wire w596;
    wire w597;
    wire w598;
    wire w599;
    wire w600;
    wire w601;
    wire w602;
    wire w603;
    wire w604;
    wire w605;
    wire w606;
    wire w607;
    wire w608;
    wire w609;
    wire w610;
    wire w611;
    wire w612;
    wire w613;
    wire w614;
    wire w615;
    wire w616;
    wire w617;
    wire w618;
    wire w619;
    wire w620;
    wire w621;
    assign out8[0] = w553;
    assign out8[1] = w554;
    assign out8[2] = w555;
    assign out8[3] = w556;
    assign out8[4] = w557;
    assign out8[5] = w558;
    assign out8[6] = w559;
    assign out8[7] = w560;
    assign out8[8] = w561;
    assign out8[9] = w562;
    assign out8[10] = w563;
    assign out8[11] = w564;
    assign out8[12] = w565;
    assign out8[13] = w566;
    assign out8[14] = w567;
    assign out8[15] = w568;
    assign out8[16] = w569;
    assign out8[17] = w570;
    assign out8[18] = w571;
    assign out8[19] = w572;
    assign out8[20] = w573;
    assign out8[21] = w574;
    assign out8[22] = w575;
    assign out8[23] = w576;
    assign out8[24] = w577;
    assign out8[25] = w578;
    assign out8[26] = w579;
    assign out8[27] = w580;
    assign out8[28] = w581;
    assign out8[29] = w582;
    assign out8[30] = w583;
    assign out8[31] = w584;
    assign out8[32] = w585;
    assign out8[33] = w586;
    assign out8[34] = w587;
    assign out8[35] = w588;
    assign out8[36] = w589;
    assign out8[37] = w590;
    assign out8[38] = w591;
    assign out8[39] = w592;
    assign out8[40] = w593;
    assign out8[41] = w594;
    assign out8[42] = w595;
    assign out8[43] = w596;
    assign out8[44] = w597;
    assign out8[45] = w598;
    assign out8[46] = w599;
    assign out8[47] = w600;
    assign out8[48] = w601;
    assign out8[49] = w602;
    assign out8[50] = w603;
    assign out8[51] = w604;
    assign out8[52] = w605;
    assign out8[53] = w606;
    assign out8[54] = w607;
    assign out8[55] = w608;
    assign out8[56] = w609;
    assign out8[57] = w610;
    assign out8[58] = w611;
    assign out8[59] = w612;
    assign out8[60] = w613;
    assign out8[61] = w614;
    assign out8[62] = w615;
    assign out8[63] = w616;
    assign out8[64] = w617;
    assign out8[65] = w618;
    assign out8[66] = w619;
    assign out8[67] = w620;
    assign out8[68] = w621;
    wire w622;
    wire w623;
    wire w624;
    wire w625;
    wire w626;
    wire w627;
    wire w628;
    wire w629;
    wire w630;
    wire w631;
    wire w632;
    wire w633;
    wire w634;
    wire w635;
    wire w636;
    wire w637;
    wire w638;
    wire w639;
    wire w640;
    wire w641;
    wire w642;
    wire w643;
    wire w644;
    wire w645;
    wire w646;
    wire w647;
    wire w648;
    wire w649;
    wire w650;
    wire w651;
    wire w652;
    wire w653;
    wire w654;
    wire w655;
    wire w656;
    wire w657;
    wire w658;
    wire w659;
    wire w660;
    wire w661;
    wire w662;
    wire w663;
    wire w664;
    wire w665;
    wire w666;
    wire w667;
    wire w668;
    wire w669;
    wire w670;
    wire w671;
    wire w672;
    wire w673;
    wire w674;
    wire w675;
    wire w676;
    wire w677;
    wire w678;
    wire w679;
    wire w680;
    wire w681;
    wire w682;
    wire w683;
    wire w684;
    wire w685;
    wire w686;
    wire w687;
    wire w688;
    wire w689;
    wire w690;
    assign out9[0] = w622;
    assign out9[1] = w623;
    assign out9[2] = w624;
    assign out9[3] = w625;
    assign out9[4] = w626;
    assign out9[5] = w627;
    assign out9[6] = w628;
    assign out9[7] = w629;
    assign out9[8] = w630;
    assign out9[9] = w631;
    assign out9[10] = w632;
    assign out9[11] = w633;
    assign out9[12] = w634;
    assign out9[13] = w635;
    assign out9[14] = w636;
    assign out9[15] = w637;
    assign out9[16] = w638;
    assign out9[17] = w639;
    assign out9[18] = w640;
    assign out9[19] = w641;
    assign out9[20] = w642;
    assign out9[21] = w643;
    assign out9[22] = w644;
    assign out9[23] = w645;
    assign out9[24] = w646;
    assign out9[25] = w647;
    assign out9[26] = w648;
    assign out9[27] = w649;
    assign out9[28] = w650;
    assign out9[29] = w651;
    assign out9[30] = w652;
    assign out9[31] = w653;
    assign out9[32] = w654;
    assign out9[33] = w655;
    assign out9[34] = w656;
    assign out9[35] = w657;
    assign out9[36] = w658;
    assign out9[37] = w659;
    assign out9[38] = w660;
    assign out9[39] = w661;
    assign out9[40] = w662;
    assign out9[41] = w663;
    assign out9[42] = w664;
    assign out9[43] = w665;
    assign out9[44] = w666;
    assign out9[45] = w667;
    assign out9[46] = w668;
    assign out9[47] = w669;
    assign out9[48] = w670;
    assign out9[49] = w671;
    assign out9[50] = w672;
    assign out9[51] = w673;
    assign out9[52] = w674;
    assign out9[53] = w675;
    assign out9[54] = w676;
    assign out9[55] = w677;
    assign out9[56] = w678;
    assign out9[57] = w679;
    assign out9[58] = w680;
    assign out9[59] = w681;
    assign out9[60] = w682;
    assign out9[61] = w683;
    assign out9[62] = w684;
    assign out9[63] = w685;
    assign out9[64] = w686;
    assign out9[65] = w687;
    assign out9[66] = w688;
    assign out9[67] = w689;
    assign out9[68] = w690;
    wire w691;
    wire w692;
    wire w693;
    wire w694;
    wire w695;
    wire w696;
    wire w697;
    wire w698;
    wire w699;
    wire w700;
    wire w701;
    wire w702;
    wire w703;
    wire w704;
    wire w705;
    wire w706;
    wire w707;
    wire w708;
    wire w709;
    wire w710;
    wire w711;
    wire w712;
    wire w713;
    wire w714;
    wire w715;
    wire w716;
    wire w717;
    wire w718;
    wire w719;
    wire w720;
    wire w721;
    wire w722;
    wire w723;
    wire w724;
    wire w725;
    wire w726;
    wire w727;
    wire w728;
    wire w729;
    wire w730;
    wire w731;
    wire w732;
    wire w733;
    wire w734;
    wire w735;
    wire w736;
    wire w737;
    wire w738;
    wire w739;
    wire w740;
    wire w741;
    wire w742;
    wire w743;
    wire w744;
    wire w745;
    wire w746;
    wire w747;
    wire w748;
    wire w749;
    wire w750;
    wire w751;
    wire w752;
    wire w753;
    wire w754;
    wire w755;
    wire w756;
    wire w757;
    wire w758;
    wire w759;
    assign out10[0] = w691;
    assign out10[1] = w692;
    assign out10[2] = w693;
    assign out10[3] = w694;
    assign out10[4] = w695;
    assign out10[5] = w696;
    assign out10[6] = w697;
    assign out10[7] = w698;
    assign out10[8] = w699;
    assign out10[9] = w700;
    assign out10[10] = w701;
    assign out10[11] = w702;
    assign out10[12] = w703;
    assign out10[13] = w704;
    assign out10[14] = w705;
    assign out10[15] = w706;
    assign out10[16] = w707;
    assign out10[17] = w708;
    assign out10[18] = w709;
    assign out10[19] = w710;
    assign out10[20] = w711;
    assign out10[21] = w712;
    assign out10[22] = w713;
    assign out10[23] = w714;
    assign out10[24] = w715;
    assign out10[25] = w716;
    assign out10[26] = w717;
    assign out10[27] = w718;
    assign out10[28] = w719;
    assign out10[29] = w720;
    assign out10[30] = w721;
    assign out10[31] = w722;
    assign out10[32] = w723;
    assign out10[33] = w724;
    assign out10[34] = w725;
    assign out10[35] = w726;
    assign out10[36] = w727;
    assign out10[37] = w728;
    assign out10[38] = w729;
    assign out10[39] = w730;
    assign out10[40] = w731;
    assign out10[41] = w732;
    assign out10[42] = w733;
    assign out10[43] = w734;
    assign out10[44] = w735;
    assign out10[45] = w736;
    assign out10[46] = w737;
    assign out10[47] = w738;
    assign out10[48] = w739;
    assign out10[49] = w740;
    assign out10[50] = w741;
    assign out10[51] = w742;
    assign out10[52] = w743;
    assign out10[53] = w744;
    assign out10[54] = w745;
    assign out10[55] = w746;
    assign out10[56] = w747;
    assign out10[57] = w748;
    assign out10[58] = w749;
    assign out10[59] = w750;
    assign out10[60] = w751;
    assign out10[61] = w752;
    assign out10[62] = w753;
    assign out10[63] = w754;
    assign out10[64] = w755;
    assign out10[65] = w756;
    assign out10[66] = w757;
    assign out10[67] = w758;
    assign out10[68] = w759;
    wire w760;
    wire w761;
    wire w762;
    wire w763;
    wire w764;
    wire w765;
    wire w766;
    wire w767;
    wire w768;
    wire w769;
    wire w770;
    wire w771;
    wire w772;
    wire w773;
    wire w774;
    wire w775;
    wire w776;
    wire w777;
    wire w778;
    wire w779;
    wire w780;
    wire w781;
    wire w782;
    wire w783;
    wire w784;
    wire w785;
    wire w786;
    wire w787;
    wire w788;
    wire w789;
    wire w790;
    wire w791;
    wire w792;
    wire w793;
    wire w794;
    wire w795;
    wire w796;
    wire w797;
    wire w798;
    wire w799;
    wire w800;
    wire w801;
    wire w802;
    wire w803;
    wire w804;
    wire w805;
    wire w806;
    wire w807;
    wire w808;
    wire w809;
    wire w810;
    wire w811;
    wire w812;
    wire w813;
    wire w814;
    wire w815;
    wire w816;
    wire w817;
    wire w818;
    wire w819;
    wire w820;
    wire w821;
    wire w822;
    wire w823;
    wire w824;
    wire w825;
    wire w826;
    wire w827;
    wire w828;
    assign out11[0] = w760;
    assign out11[1] = w761;
    assign out11[2] = w762;
    assign out11[3] = w763;
    assign out11[4] = w764;
    assign out11[5] = w765;
    assign out11[6] = w766;
    assign out11[7] = w767;
    assign out11[8] = w768;
    assign out11[9] = w769;
    assign out11[10] = w770;
    assign out11[11] = w771;
    assign out11[12] = w772;
    assign out11[13] = w773;
    assign out11[14] = w774;
    assign out11[15] = w775;
    assign out11[16] = w776;
    assign out11[17] = w777;
    assign out11[18] = w778;
    assign out11[19] = w779;
    assign out11[20] = w780;
    assign out11[21] = w781;
    assign out11[22] = w782;
    assign out11[23] = w783;
    assign out11[24] = w784;
    assign out11[25] = w785;
    assign out11[26] = w786;
    assign out11[27] = w787;
    assign out11[28] = w788;
    assign out11[29] = w789;
    assign out11[30] = w790;
    assign out11[31] = w791;
    assign out11[32] = w792;
    assign out11[33] = w793;
    assign out11[34] = w794;
    assign out11[35] = w795;
    assign out11[36] = w796;
    assign out11[37] = w797;
    assign out11[38] = w798;
    assign out11[39] = w799;
    assign out11[40] = w800;
    assign out11[41] = w801;
    assign out11[42] = w802;
    assign out11[43] = w803;
    assign out11[44] = w804;
    assign out11[45] = w805;
    assign out11[46] = w806;
    assign out11[47] = w807;
    assign out11[48] = w808;
    assign out11[49] = w809;
    assign out11[50] = w810;
    assign out11[51] = w811;
    assign out11[52] = w812;
    assign out11[53] = w813;
    assign out11[54] = w814;
    assign out11[55] = w815;
    assign out11[56] = w816;
    assign out11[57] = w817;
    assign out11[58] = w818;
    assign out11[59] = w819;
    assign out11[60] = w820;
    assign out11[61] = w821;
    assign out11[62] = w822;
    assign out11[63] = w823;
    assign out11[64] = w824;
    assign out11[65] = w825;
    assign out11[66] = w826;
    assign out11[67] = w827;
    assign out11[68] = w828;
    wire w829;
    wire w830;
    wire w831;
    wire w832;
    wire w833;
    wire w834;
    wire w835;
    wire w836;
    wire w837;
    wire w838;
    wire w839;
    wire w840;
    wire w841;
    wire w842;
    wire w843;
    wire w844;
    wire w845;
    wire w846;
    wire w847;
    wire w848;
    wire w849;
    wire w850;
    wire w851;
    wire w852;
    wire w853;
    wire w854;
    wire w855;
    wire w856;
    wire w857;
    wire w858;
    wire w859;
    wire w860;
    wire w861;
    wire w862;
    wire w863;
    wire w864;
    wire w865;
    wire w866;
    wire w867;
    wire w868;
    wire w869;
    wire w870;
    wire w871;
    wire w872;
    wire w873;
    wire w874;
    wire w875;
    wire w876;
    wire w877;
    wire w878;
    wire w879;
    wire w880;
    wire w881;
    wire w882;
    wire w883;
    wire w884;
    wire w885;
    wire w886;
    wire w887;
    wire w888;
    wire w889;
    wire w890;
    wire w891;
    wire w892;
    wire w893;
    wire w894;
    wire w895;
    wire w896;
    wire w897;
    assign out12[0] = w829;
    assign out12[1] = w830;
    assign out12[2] = w831;
    assign out12[3] = w832;
    assign out12[4] = w833;
    assign out12[5] = w834;
    assign out12[6] = w835;
    assign out12[7] = w836;
    assign out12[8] = w837;
    assign out12[9] = w838;
    assign out12[10] = w839;
    assign out12[11] = w840;
    assign out12[12] = w841;
    assign out12[13] = w842;
    assign out12[14] = w843;
    assign out12[15] = w844;
    assign out12[16] = w845;
    assign out12[17] = w846;
    assign out12[18] = w847;
    assign out12[19] = w848;
    assign out12[20] = w849;
    assign out12[21] = w850;
    assign out12[22] = w851;
    assign out12[23] = w852;
    assign out12[24] = w853;
    assign out12[25] = w854;
    assign out12[26] = w855;
    assign out12[27] = w856;
    assign out12[28] = w857;
    assign out12[29] = w858;
    assign out12[30] = w859;
    assign out12[31] = w860;
    assign out12[32] = w861;
    assign out12[33] = w862;
    assign out12[34] = w863;
    assign out12[35] = w864;
    assign out12[36] = w865;
    assign out12[37] = w866;
    assign out12[38] = w867;
    assign out12[39] = w868;
    assign out12[40] = w869;
    assign out12[41] = w870;
    assign out12[42] = w871;
    assign out12[43] = w872;
    assign out12[44] = w873;
    assign out12[45] = w874;
    assign out12[46] = w875;
    assign out12[47] = w876;
    assign out12[48] = w877;
    assign out12[49] = w878;
    assign out12[50] = w879;
    assign out12[51] = w880;
    assign out12[52] = w881;
    assign out12[53] = w882;
    assign out12[54] = w883;
    assign out12[55] = w884;
    assign out12[56] = w885;
    assign out12[57] = w886;
    assign out12[58] = w887;
    assign out12[59] = w888;
    assign out12[60] = w889;
    assign out12[61] = w890;
    assign out12[62] = w891;
    assign out12[63] = w892;
    assign out12[64] = w893;
    assign out12[65] = w894;
    assign out12[66] = w895;
    assign out12[67] = w896;
    assign out12[68] = w897;
    wire w898;
    wire w899;
    wire w900;
    wire w901;
    wire w902;
    wire w903;
    wire w904;
    wire w905;
    wire w906;
    wire w907;
    wire w908;
    wire w909;
    wire w910;
    wire w911;
    wire w912;
    wire w913;
    wire w914;
    wire w915;
    wire w916;
    wire w917;
    wire w918;
    wire w919;
    wire w920;
    wire w921;
    wire w922;
    wire w923;
    wire w924;
    wire w925;
    wire w926;
    wire w927;
    wire w928;
    wire w929;
    wire w930;
    wire w931;
    wire w932;
    wire w933;
    wire w934;
    wire w935;
    wire w936;
    wire w937;
    wire w938;
    wire w939;
    wire w940;
    wire w941;
    wire w942;
    wire w943;
    wire w944;
    wire w945;
    wire w946;
    wire w947;
    wire w948;
    wire w949;
    wire w950;
    wire w951;
    wire w952;
    wire w953;
    wire w954;
    wire w955;
    wire w956;
    wire w957;
    wire w958;
    wire w959;
    wire w960;
    wire w961;
    wire w962;
    wire w963;
    wire w964;
    wire w965;
    wire w966;
    assign out13[0] = w898;
    assign out13[1] = w899;
    assign out13[2] = w900;
    assign out13[3] = w901;
    assign out13[4] = w902;
    assign out13[5] = w903;
    assign out13[6] = w904;
    assign out13[7] = w905;
    assign out13[8] = w906;
    assign out13[9] = w907;
    assign out13[10] = w908;
    assign out13[11] = w909;
    assign out13[12] = w910;
    assign out13[13] = w911;
    assign out13[14] = w912;
    assign out13[15] = w913;
    assign out13[16] = w914;
    assign out13[17] = w915;
    assign out13[18] = w916;
    assign out13[19] = w917;
    assign out13[20] = w918;
    assign out13[21] = w919;
    assign out13[22] = w920;
    assign out13[23] = w921;
    assign out13[24] = w922;
    assign out13[25] = w923;
    assign out13[26] = w924;
    assign out13[27] = w925;
    assign out13[28] = w926;
    assign out13[29] = w927;
    assign out13[30] = w928;
    assign out13[31] = w929;
    assign out13[32] = w930;
    assign out13[33] = w931;
    assign out13[34] = w932;
    assign out13[35] = w933;
    assign out13[36] = w934;
    assign out13[37] = w935;
    assign out13[38] = w936;
    assign out13[39] = w937;
    assign out13[40] = w938;
    assign out13[41] = w939;
    assign out13[42] = w940;
    assign out13[43] = w941;
    assign out13[44] = w942;
    assign out13[45] = w943;
    assign out13[46] = w944;
    assign out13[47] = w945;
    assign out13[48] = w946;
    assign out13[49] = w947;
    assign out13[50] = w948;
    assign out13[51] = w949;
    assign out13[52] = w950;
    assign out13[53] = w951;
    assign out13[54] = w952;
    assign out13[55] = w953;
    assign out13[56] = w954;
    assign out13[57] = w955;
    assign out13[58] = w956;
    assign out13[59] = w957;
    assign out13[60] = w958;
    assign out13[61] = w959;
    assign out13[62] = w960;
    assign out13[63] = w961;
    assign out13[64] = w962;
    assign out13[65] = w963;
    assign out13[66] = w964;
    assign out13[67] = w965;
    assign out13[68] = w966;
    wire w967;
    wire w968;
    wire w969;
    wire w970;
    wire w971;
    wire w972;
    wire w973;
    wire w974;
    wire w975;
    wire w976;
    wire w977;
    wire w978;
    wire w979;
    wire w980;
    wire w981;
    wire w982;
    wire w983;
    wire w984;
    wire w985;
    wire w986;
    wire w987;
    wire w988;
    wire w989;
    wire w990;
    wire w991;
    wire w992;
    wire w993;
    wire w994;
    wire w995;
    wire w996;
    wire w997;
    wire w998;
    wire w999;
    wire w1000;
    wire w1001;
    wire w1002;
    wire w1003;
    wire w1004;
    wire w1005;
    wire w1006;
    wire w1007;
    wire w1008;
    wire w1009;
    wire w1010;
    wire w1011;
    wire w1012;
    wire w1013;
    wire w1014;
    wire w1015;
    wire w1016;
    wire w1017;
    wire w1018;
    wire w1019;
    wire w1020;
    wire w1021;
    wire w1022;
    wire w1023;
    wire w1024;
    wire w1025;
    wire w1026;
    wire w1027;
    wire w1028;
    wire w1029;
    wire w1030;
    wire w1031;
    wire w1032;
    wire w1033;
    wire w1034;
    wire w1035;
    assign out14[0] = w967;
    assign out14[1] = w968;
    assign out14[2] = w969;
    assign out14[3] = w970;
    assign out14[4] = w971;
    assign out14[5] = w972;
    assign out14[6] = w973;
    assign out14[7] = w974;
    assign out14[8] = w975;
    assign out14[9] = w976;
    assign out14[10] = w977;
    assign out14[11] = w978;
    assign out14[12] = w979;
    assign out14[13] = w980;
    assign out14[14] = w981;
    assign out14[15] = w982;
    assign out14[16] = w983;
    assign out14[17] = w984;
    assign out14[18] = w985;
    assign out14[19] = w986;
    assign out14[20] = w987;
    assign out14[21] = w988;
    assign out14[22] = w989;
    assign out14[23] = w990;
    assign out14[24] = w991;
    assign out14[25] = w992;
    assign out14[26] = w993;
    assign out14[27] = w994;
    assign out14[28] = w995;
    assign out14[29] = w996;
    assign out14[30] = w997;
    assign out14[31] = w998;
    assign out14[32] = w999;
    assign out14[33] = w1000;
    assign out14[34] = w1001;
    assign out14[35] = w1002;
    assign out14[36] = w1003;
    assign out14[37] = w1004;
    assign out14[38] = w1005;
    assign out14[39] = w1006;
    assign out14[40] = w1007;
    assign out14[41] = w1008;
    assign out14[42] = w1009;
    assign out14[43] = w1010;
    assign out14[44] = w1011;
    assign out14[45] = w1012;
    assign out14[46] = w1013;
    assign out14[47] = w1014;
    assign out14[48] = w1015;
    assign out14[49] = w1016;
    assign out14[50] = w1017;
    assign out14[51] = w1018;
    assign out14[52] = w1019;
    assign out14[53] = w1020;
    assign out14[54] = w1021;
    assign out14[55] = w1022;
    assign out14[56] = w1023;
    assign out14[57] = w1024;
    assign out14[58] = w1025;
    assign out14[59] = w1026;
    assign out14[60] = w1027;
    assign out14[61] = w1028;
    assign out14[62] = w1029;
    assign out14[63] = w1030;
    assign out14[64] = w1031;
    assign out14[65] = w1032;
    assign out14[66] = w1033;
    assign out14[67] = w1034;
    assign out14[68] = w1035;
    wire w1036;
    wire w1037;
    wire w1038;
    wire w1039;
    wire w1040;
    wire w1041;
    wire w1042;
    wire w1043;
    wire w1044;
    wire w1045;
    wire w1046;
    wire w1047;
    wire w1048;
    wire w1049;
    wire w1050;
    wire w1051;
    wire w1052;
    wire w1053;
    wire w1054;
    wire w1055;
    wire w1056;
    wire w1057;
    wire w1058;
    wire w1059;
    wire w1060;
    wire w1061;
    wire w1062;
    wire w1063;
    wire w1064;
    wire w1065;
    wire w1066;
    wire w1067;
    wire w1068;
    wire w1069;
    wire w1070;
    wire w1071;
    wire w1072;
    wire w1073;
    wire w1074;
    wire w1075;
    wire w1076;
    wire w1077;
    wire w1078;
    wire w1079;
    wire w1080;
    wire w1081;
    wire w1082;
    wire w1083;
    wire w1084;
    wire w1085;
    wire w1086;
    wire w1087;
    wire w1088;
    wire w1089;
    wire w1090;
    wire w1091;
    wire w1092;
    wire w1093;
    wire w1094;
    wire w1095;
    wire w1096;
    wire w1097;
    wire w1098;
    wire w1099;
    wire w1100;
    wire w1101;
    wire w1102;
    wire w1103;
    wire w1104;
    assign out15[0] = w1036;
    assign out15[1] = w1037;
    assign out15[2] = w1038;
    assign out15[3] = w1039;
    assign out15[4] = w1040;
    assign out15[5] = w1041;
    assign out15[6] = w1042;
    assign out15[7] = w1043;
    assign out15[8] = w1044;
    assign out15[9] = w1045;
    assign out15[10] = w1046;
    assign out15[11] = w1047;
    assign out15[12] = w1048;
    assign out15[13] = w1049;
    assign out15[14] = w1050;
    assign out15[15] = w1051;
    assign out15[16] = w1052;
    assign out15[17] = w1053;
    assign out15[18] = w1054;
    assign out15[19] = w1055;
    assign out15[20] = w1056;
    assign out15[21] = w1057;
    assign out15[22] = w1058;
    assign out15[23] = w1059;
    assign out15[24] = w1060;
    assign out15[25] = w1061;
    assign out15[26] = w1062;
    assign out15[27] = w1063;
    assign out15[28] = w1064;
    assign out15[29] = w1065;
    assign out15[30] = w1066;
    assign out15[31] = w1067;
    assign out15[32] = w1068;
    assign out15[33] = w1069;
    assign out15[34] = w1070;
    assign out15[35] = w1071;
    assign out15[36] = w1072;
    assign out15[37] = w1073;
    assign out15[38] = w1074;
    assign out15[39] = w1075;
    assign out15[40] = w1076;
    assign out15[41] = w1077;
    assign out15[42] = w1078;
    assign out15[43] = w1079;
    assign out15[44] = w1080;
    assign out15[45] = w1081;
    assign out15[46] = w1082;
    assign out15[47] = w1083;
    assign out15[48] = w1084;
    assign out15[49] = w1085;
    assign out15[50] = w1086;
    assign out15[51] = w1087;
    assign out15[52] = w1088;
    assign out15[53] = w1089;
    assign out15[54] = w1090;
    assign out15[55] = w1091;
    assign out15[56] = w1092;
    assign out15[57] = w1093;
    assign out15[58] = w1094;
    assign out15[59] = w1095;
    assign out15[60] = w1096;
    assign out15[61] = w1097;
    assign out15[62] = w1098;
    assign out15[63] = w1099;
    assign out15[64] = w1100;
    assign out15[65] = w1101;
    assign out15[66] = w1102;
    assign out15[67] = w1103;
    assign out15[68] = w1104;
    sw_m #(.SIZE(69)) sw0({w69,w68,w67,w66,w65,w64,w63,w62,w61,w60,w59,w58,w57,w56,w55,w54,w53,w52,w51,w50,w49,w48,w47,w46,w45,w44,w43,w42,w41,w40,w39,w38,w37,w36,w35,w34,w33,w32,w31,w30,w29,w28,w27,w26,w25,w24,w23,w22,w21,w20,w19,w18,w17,w16,w15,w14,w13,w12,w11,w10,w9,w8,w7,w6,w5,w4,w3,w2,w1}, {w138,w137,w136,w135,w134,w133,w132,w131,w130,w129,w128,w127,w126,w125,w124,w123,w122,w121,w120,w119,w118,w117,w116,w115,w114,w113,w112,w111,w110,w109,w108,w107,w106,w105,w104,w103,w102,w101,w100,w99,w98,w97,w96,w95,w94,w93,w92,w91,w90,w89,w88,w87,w86,w85,w84,w83,w82,w81,w80,w79,w78,w77,w76,w75,w74,w73,w72,w71,w70}, x0_69, {x0_68,x0_67,x0_66,x0_65,x0_64,x0_63,x0_62,x0_61,x0_60,x0_59,x0_58,x0_57,x0_56,x0_55,x0_54,x0_53,x0_52,x0_51,x0_50,x0_49,x0_48,x0_47,x0_46,x0_45,x0_44,x0_43,x0_42,x0_41,x0_40,x0_39,x0_38,x0_37,x0_36,x0_35,x0_34,x0_33,x0_32,x0_31,x0_30,x0_29,x0_28,x0_27,x0_26,x0_25,x0_24,x0_23,x0_22,x0_21,x0_20,x0_19,x0_18,x0_17,x0_16,x0_15,x0_14,x0_13,x0_12,x0_11,x0_10,x0_9,x0_8,x0_7,x0_6,x0_5,x0_4,x0_3,x0_2,x0_1,x0_0}, {x1_68,x1_67,x1_66,x1_65,x1_64,x1_63,x1_62,x1_61,x1_60,x1_59,x1_58,x1_57,x1_56,x1_55,x1_54,x1_53,x1_52,x1_51,x1_50,x1_49,x1_48,x1_47,x1_46,x1_45,x1_44,x1_43,x1_42,x1_41,x1_40,x1_39,x1_38,x1_37,x1_36,x1_35,x1_34,x1_33,x1_32,x1_31,x1_30,x1_29,x1_28,x1_27,x1_26,x1_25,x1_24,x1_23,x1_22,x1_21,x1_20,x1_19,x1_18,x1_17,x1_16,x1_15,x1_14,x1_13,x1_12,x1_11,x1_10,x1_9,x1_8,x1_7,x1_6,x1_5,x1_4,x1_3,x1_2,x1_1,x1_0});
    sw_m #(.SIZE(69)) sw1({w759,w758,w757,w756,w755,w754,w753,w752,w751,w750,w749,w748,w747,w746,w745,w744,w743,w742,w741,w740,w739,w738,w737,w736,w735,w734,w733,w732,w731,w730,w729,w728,w727,w726,w725,w724,w723,w722,w721,w720,w719,w718,w717,w716,w715,w714,w713,w712,w711,w710,w709,w708,w707,w706,w705,w704,w703,w702,w701,w700,w699,w698,w697,w696,w695,w694,w693,w692,w691}, {w828,w827,w826,w825,w824,w823,w822,w821,w820,w819,w818,w817,w816,w815,w814,w813,w812,w811,w810,w809,w808,w807,w806,w805,w804,w803,w802,w801,w800,w799,w798,w797,w796,w795,w794,w793,w792,w791,w790,w789,w788,w787,w786,w785,w784,w783,w782,w781,w780,w779,w778,w777,w776,w775,w774,w773,w772,w771,w770,w769,w768,w767,w766,w765,w764,w763,w762,w761,w760}, x10_69, {x10_68,x10_67,x10_66,x10_65,x10_64,x10_63,x10_62,x10_61,x10_60,x10_59,x10_58,x10_57,x10_56,x10_55,x10_54,x10_53,x10_52,x10_51,x10_50,x10_49,x10_48,x10_47,x10_46,x10_45,x10_44,x10_43,x10_42,x10_41,x10_40,x10_39,x10_38,x10_37,x10_36,x10_35,x10_34,x10_33,x10_32,x10_31,x10_30,x10_29,x10_28,x10_27,x10_26,x10_25,x10_24,x10_23,x10_22,x10_21,x10_20,x10_19,x10_18,x10_17,x10_16,x10_15,x10_14,x10_13,x10_12,x10_11,x10_10,x10_9,x10_8,x10_7,x10_6,x10_5,x10_4,x10_3,x10_2,x10_1,x10_0}, {x11_68,x11_67,x11_66,x11_65,x11_64,x11_63,x11_62,x11_61,x11_60,x11_59,x11_58,x11_57,x11_56,x11_55,x11_54,x11_53,x11_52,x11_51,x11_50,x11_49,x11_48,x11_47,x11_46,x11_45,x11_44,x11_43,x11_42,x11_41,x11_40,x11_39,x11_38,x11_37,x11_36,x11_35,x11_34,x11_33,x11_32,x11_31,x11_30,x11_29,x11_28,x11_27,x11_26,x11_25,x11_24,x11_23,x11_22,x11_21,x11_20,x11_19,x11_18,x11_17,x11_16,x11_15,x11_14,x11_13,x11_12,x11_11,x11_10,x11_9,x11_8,x11_7,x11_6,x11_5,x11_4,x11_3,x11_2,x11_1,x11_0});
    sw_m #(.SIZE(69)) sw2({w897,w896,w895,w894,w893,w892,w891,w890,w889,w888,w887,w886,w885,w884,w883,w882,w881,w880,w879,w878,w877,w876,w875,w874,w873,w872,w871,w870,w869,w868,w867,w866,w865,w864,w863,w862,w861,w860,w859,w858,w857,w856,w855,w854,w853,w852,w851,w850,w849,w848,w847,w846,w845,w844,w843,w842,w841,w840,w839,w838,w837,w836,w835,w834,w833,w832,w831,w830,w829}, {w966,w965,w964,w963,w962,w961,w960,w959,w958,w957,w956,w955,w954,w953,w952,w951,w950,w949,w948,w947,w946,w945,w944,w943,w942,w941,w940,w939,w938,w937,w936,w935,w934,w933,w932,w931,w930,w929,w928,w927,w926,w925,w924,w923,w922,w921,w920,w919,w918,w917,w916,w915,w914,w913,w912,w911,w910,w909,w908,w907,w906,w905,w904,w903,w902,w901,w900,w899,w898}, x12_69, {x12_68,x12_67,x12_66,x12_65,x12_64,x12_63,x12_62,x12_61,x12_60,x12_59,x12_58,x12_57,x12_56,x12_55,x12_54,x12_53,x12_52,x12_51,x12_50,x12_49,x12_48,x12_47,x12_46,x12_45,x12_44,x12_43,x12_42,x12_41,x12_40,x12_39,x12_38,x12_37,x12_36,x12_35,x12_34,x12_33,x12_32,x12_31,x12_30,x12_29,x12_28,x12_27,x12_26,x12_25,x12_24,x12_23,x12_22,x12_21,x12_20,x12_19,x12_18,x12_17,x12_16,x12_15,x12_14,x12_13,x12_12,x12_11,x12_10,x12_9,x12_8,x12_7,x12_6,x12_5,x12_4,x12_3,x12_2,x12_1,x12_0}, {x13_68,x13_67,x13_66,x13_65,x13_64,x13_63,x13_62,x13_61,x13_60,x13_59,x13_58,x13_57,x13_56,x13_55,x13_54,x13_53,x13_52,x13_51,x13_50,x13_49,x13_48,x13_47,x13_46,x13_45,x13_44,x13_43,x13_42,x13_41,x13_40,x13_39,x13_38,x13_37,x13_36,x13_35,x13_34,x13_33,x13_32,x13_31,x13_30,x13_29,x13_28,x13_27,x13_26,x13_25,x13_24,x13_23,x13_22,x13_21,x13_20,x13_19,x13_18,x13_17,x13_16,x13_15,x13_14,x13_13,x13_12,x13_11,x13_10,x13_9,x13_8,x13_7,x13_6,x13_5,x13_4,x13_3,x13_2,x13_1,x13_0});
    sw_m #(.SIZE(69)) sw3({w1035,w1034,w1033,w1032,w1031,w1030,w1029,w1028,w1027,w1026,w1025,w1024,w1023,w1022,w1021,w1020,w1019,w1018,w1017,w1016,w1015,w1014,w1013,w1012,w1011,w1010,w1009,w1008,w1007,w1006,w1005,w1004,w1003,w1002,w1001,w1000,w999,w998,w997,w996,w995,w994,w993,w992,w991,w990,w989,w988,w987,w986,w985,w984,w983,w982,w981,w980,w979,w978,w977,w976,w975,w974,w973,w972,w971,w970,w969,w968,w967}, {w1104,w1103,w1102,w1101,w1100,w1099,w1098,w1097,w1096,w1095,w1094,w1093,w1092,w1091,w1090,w1089,w1088,w1087,w1086,w1085,w1084,w1083,w1082,w1081,w1080,w1079,w1078,w1077,w1076,w1075,w1074,w1073,w1072,w1071,w1070,w1069,w1068,w1067,w1066,w1065,w1064,w1063,w1062,w1061,w1060,w1059,w1058,w1057,w1056,w1055,w1054,w1053,w1052,w1051,w1050,w1049,w1048,w1047,w1046,w1045,w1044,w1043,w1042,w1041,w1040,w1039,w1038,w1037,w1036}, x14_69, {x14_68,x14_67,x14_66,x14_65,x14_64,x14_63,x14_62,x14_61,x14_60,x14_59,x14_58,x14_57,x14_56,x14_55,x14_54,x14_53,x14_52,x14_51,x14_50,x14_49,x14_48,x14_47,x14_46,x14_45,x14_44,x14_43,x14_42,x14_41,x14_40,x14_39,x14_38,x14_37,x14_36,x14_35,x14_34,x14_33,x14_32,x14_31,x14_30,x14_29,x14_28,x14_27,x14_26,x14_25,x14_24,x14_23,x14_22,x14_21,x14_20,x14_19,x14_18,x14_17,x14_16,x14_15,x14_14,x14_13,x14_12,x14_11,x14_10,x14_9,x14_8,x14_7,x14_6,x14_5,x14_4,x14_3,x14_2,x14_1,x14_0}, {x15_68,x15_67,x15_66,x15_65,x15_64,x15_63,x15_62,x15_61,x15_60,x15_59,x15_58,x15_57,x15_56,x15_55,x15_54,x15_53,x15_52,x15_51,x15_50,x15_49,x15_48,x15_47,x15_46,x15_45,x15_44,x15_43,x15_42,x15_41,x15_40,x15_39,x15_38,x15_37,x15_36,x15_35,x15_34,x15_33,x15_32,x15_31,x15_30,x15_29,x15_28,x15_27,x15_26,x15_25,x15_24,x15_23,x15_22,x15_21,x15_20,x15_19,x15_18,x15_17,x15_16,x15_15,x15_14,x15_13,x15_12,x15_11,x15_10,x15_9,x15_8,x15_7,x15_6,x15_5,x15_4,x15_3,x15_2,x15_1,x15_0});
    sw_m #(.SIZE(69)) sw4({w207,w206,w205,w204,w203,w202,w201,w200,w199,w198,w197,w196,w195,w194,w193,w192,w191,w190,w189,w188,w187,w186,w185,w184,w183,w182,w181,w180,w179,w178,w177,w176,w175,w174,w173,w172,w171,w170,w169,w168,w167,w166,w165,w164,w163,w162,w161,w160,w159,w158,w157,w156,w155,w154,w153,w152,w151,w150,w149,w148,w147,w146,w145,w144,w143,w142,w141,w140,w139}, {w276,w275,w274,w273,w272,w271,w270,w269,w268,w267,w266,w265,w264,w263,w262,w261,w260,w259,w258,w257,w256,w255,w254,w253,w252,w251,w250,w249,w248,w247,w246,w245,w244,w243,w242,w241,w240,w239,w238,w237,w236,w235,w234,w233,w232,w231,w230,w229,w228,w227,w226,w225,w224,w223,w222,w221,w220,w219,w218,w217,w216,w215,w214,w213,w212,w211,w210,w209,w208}, x2_69, {x2_68,x2_67,x2_66,x2_65,x2_64,x2_63,x2_62,x2_61,x2_60,x2_59,x2_58,x2_57,x2_56,x2_55,x2_54,x2_53,x2_52,x2_51,x2_50,x2_49,x2_48,x2_47,x2_46,x2_45,x2_44,x2_43,x2_42,x2_41,x2_40,x2_39,x2_38,x2_37,x2_36,x2_35,x2_34,x2_33,x2_32,x2_31,x2_30,x2_29,x2_28,x2_27,x2_26,x2_25,x2_24,x2_23,x2_22,x2_21,x2_20,x2_19,x2_18,x2_17,x2_16,x2_15,x2_14,x2_13,x2_12,x2_11,x2_10,x2_9,x2_8,x2_7,x2_6,x2_5,x2_4,x2_3,x2_2,x2_1,x2_0}, {x3_68,x3_67,x3_66,x3_65,x3_64,x3_63,x3_62,x3_61,x3_60,x3_59,x3_58,x3_57,x3_56,x3_55,x3_54,x3_53,x3_52,x3_51,x3_50,x3_49,x3_48,x3_47,x3_46,x3_45,x3_44,x3_43,x3_42,x3_41,x3_40,x3_39,x3_38,x3_37,x3_36,x3_35,x3_34,x3_33,x3_32,x3_31,x3_30,x3_29,x3_28,x3_27,x3_26,x3_25,x3_24,x3_23,x3_22,x3_21,x3_20,x3_19,x3_18,x3_17,x3_16,x3_15,x3_14,x3_13,x3_12,x3_11,x3_10,x3_9,x3_8,x3_7,x3_6,x3_5,x3_4,x3_3,x3_2,x3_1,x3_0});
    sw_m #(.SIZE(69)) sw5({w345,w344,w343,w342,w341,w340,w339,w338,w337,w336,w335,w334,w333,w332,w331,w330,w329,w328,w327,w326,w325,w324,w323,w322,w321,w320,w319,w318,w317,w316,w315,w314,w313,w312,w311,w310,w309,w308,w307,w306,w305,w304,w303,w302,w301,w300,w299,w298,w297,w296,w295,w294,w293,w292,w291,w290,w289,w288,w287,w286,w285,w284,w283,w282,w281,w280,w279,w278,w277}, {w414,w413,w412,w411,w410,w409,w408,w407,w406,w405,w404,w403,w402,w401,w400,w399,w398,w397,w396,w395,w394,w393,w392,w391,w390,w389,w388,w387,w386,w385,w384,w383,w382,w381,w380,w379,w378,w377,w376,w375,w374,w373,w372,w371,w370,w369,w368,w367,w366,w365,w364,w363,w362,w361,w360,w359,w358,w357,w356,w355,w354,w353,w352,w351,w350,w349,w348,w347,w346}, x4_69, {x4_68,x4_67,x4_66,x4_65,x4_64,x4_63,x4_62,x4_61,x4_60,x4_59,x4_58,x4_57,x4_56,x4_55,x4_54,x4_53,x4_52,x4_51,x4_50,x4_49,x4_48,x4_47,x4_46,x4_45,x4_44,x4_43,x4_42,x4_41,x4_40,x4_39,x4_38,x4_37,x4_36,x4_35,x4_34,x4_33,x4_32,x4_31,x4_30,x4_29,x4_28,x4_27,x4_26,x4_25,x4_24,x4_23,x4_22,x4_21,x4_20,x4_19,x4_18,x4_17,x4_16,x4_15,x4_14,x4_13,x4_12,x4_11,x4_10,x4_9,x4_8,x4_7,x4_6,x4_5,x4_4,x4_3,x4_2,x4_1,x4_0}, {x5_68,x5_67,x5_66,x5_65,x5_64,x5_63,x5_62,x5_61,x5_60,x5_59,x5_58,x5_57,x5_56,x5_55,x5_54,x5_53,x5_52,x5_51,x5_50,x5_49,x5_48,x5_47,x5_46,x5_45,x5_44,x5_43,x5_42,x5_41,x5_40,x5_39,x5_38,x5_37,x5_36,x5_35,x5_34,x5_33,x5_32,x5_31,x5_30,x5_29,x5_28,x5_27,x5_26,x5_25,x5_24,x5_23,x5_22,x5_21,x5_20,x5_19,x5_18,x5_17,x5_16,x5_15,x5_14,x5_13,x5_12,x5_11,x5_10,x5_9,x5_8,x5_7,x5_6,x5_5,x5_4,x5_3,x5_2,x5_1,x5_0});
    sw_m #(.SIZE(69)) sw6({w483,w482,w481,w480,w479,w478,w477,w476,w475,w474,w473,w472,w471,w470,w469,w468,w467,w466,w465,w464,w463,w462,w461,w460,w459,w458,w457,w456,w455,w454,w453,w452,w451,w450,w449,w448,w447,w446,w445,w444,w443,w442,w441,w440,w439,w438,w437,w436,w435,w434,w433,w432,w431,w430,w429,w428,w427,w426,w425,w424,w423,w422,w421,w420,w419,w418,w417,w416,w415}, {w552,w551,w550,w549,w548,w547,w546,w545,w544,w543,w542,w541,w540,w539,w538,w537,w536,w535,w534,w533,w532,w531,w530,w529,w528,w527,w526,w525,w524,w523,w522,w521,w520,w519,w518,w517,w516,w515,w514,w513,w512,w511,w510,w509,w508,w507,w506,w505,w504,w503,w502,w501,w500,w499,w498,w497,w496,w495,w494,w493,w492,w491,w490,w489,w488,w487,w486,w485,w484}, x6_69, {x6_68,x6_67,x6_66,x6_65,x6_64,x6_63,x6_62,x6_61,x6_60,x6_59,x6_58,x6_57,x6_56,x6_55,x6_54,x6_53,x6_52,x6_51,x6_50,x6_49,x6_48,x6_47,x6_46,x6_45,x6_44,x6_43,x6_42,x6_41,x6_40,x6_39,x6_38,x6_37,x6_36,x6_35,x6_34,x6_33,x6_32,x6_31,x6_30,x6_29,x6_28,x6_27,x6_26,x6_25,x6_24,x6_23,x6_22,x6_21,x6_20,x6_19,x6_18,x6_17,x6_16,x6_15,x6_14,x6_13,x6_12,x6_11,x6_10,x6_9,x6_8,x6_7,x6_6,x6_5,x6_4,x6_3,x6_2,x6_1,x6_0}, {x7_68,x7_67,x7_66,x7_65,x7_64,x7_63,x7_62,x7_61,x7_60,x7_59,x7_58,x7_57,x7_56,x7_55,x7_54,x7_53,x7_52,x7_51,x7_50,x7_49,x7_48,x7_47,x7_46,x7_45,x7_44,x7_43,x7_42,x7_41,x7_40,x7_39,x7_38,x7_37,x7_36,x7_35,x7_34,x7_33,x7_32,x7_31,x7_30,x7_29,x7_28,x7_27,x7_26,x7_25,x7_24,x7_23,x7_22,x7_21,x7_20,x7_19,x7_18,x7_17,x7_16,x7_15,x7_14,x7_13,x7_12,x7_11,x7_10,x7_9,x7_8,x7_7,x7_6,x7_5,x7_4,x7_3,x7_2,x7_1,x7_0});
    sw_m #(.SIZE(69)) sw7({w621,w620,w619,w618,w617,w616,w615,w614,w613,w612,w611,w610,w609,w608,w607,w606,w605,w604,w603,w602,w601,w600,w599,w598,w597,w596,w595,w594,w593,w592,w591,w590,w589,w588,w587,w586,w585,w584,w583,w582,w581,w580,w579,w578,w577,w576,w575,w574,w573,w572,w571,w570,w569,w568,w567,w566,w565,w564,w563,w562,w561,w560,w559,w558,w557,w556,w555,w554,w553}, {w690,w689,w688,w687,w686,w685,w684,w683,w682,w681,w680,w679,w678,w677,w676,w675,w674,w673,w672,w671,w670,w669,w668,w667,w666,w665,w664,w663,w662,w661,w660,w659,w658,w657,w656,w655,w654,w653,w652,w651,w650,w649,w648,w647,w646,w645,w644,w643,w642,w641,w640,w639,w638,w637,w636,w635,w634,w633,w632,w631,w630,w629,w628,w627,w626,w625,w624,w623,w622}, x8_69, {x8_68,x8_67,x8_66,x8_65,x8_64,x8_63,x8_62,x8_61,x8_60,x8_59,x8_58,x8_57,x8_56,x8_55,x8_54,x8_53,x8_52,x8_51,x8_50,x8_49,x8_48,x8_47,x8_46,x8_45,x8_44,x8_43,x8_42,x8_41,x8_40,x8_39,x8_38,x8_37,x8_36,x8_35,x8_34,x8_33,x8_32,x8_31,x8_30,x8_29,x8_28,x8_27,x8_26,x8_25,x8_24,x8_23,x8_22,x8_21,x8_20,x8_19,x8_18,x8_17,x8_16,x8_15,x8_14,x8_13,x8_12,x8_11,x8_10,x8_9,x8_8,x8_7,x8_6,x8_5,x8_4,x8_3,x8_2,x8_1,x8_0}, {x9_68,x9_67,x9_66,x9_65,x9_64,x9_63,x9_62,x9_61,x9_60,x9_59,x9_58,x9_57,x9_56,x9_55,x9_54,x9_53,x9_52,x9_51,x9_50,x9_49,x9_48,x9_47,x9_46,x9_45,x9_44,x9_43,x9_42,x9_41,x9_40,x9_39,x9_38,x9_37,x9_36,x9_35,x9_34,x9_33,x9_32,x9_31,x9_30,x9_29,x9_28,x9_27,x9_26,x9_25,x9_24,x9_23,x9_22,x9_21,x9_20,x9_19,x9_18,x9_17,x9_16,x9_15,x9_14,x9_13,x9_12,x9_11,x9_10,x9_9,x9_8,x9_7,x9_6,x9_5,x9_4,x9_3,x9_2,x9_1,x9_0});
endmodule
