`default_nettype none

module parPrefix2OR_16 (
output wire [16-1:0] out,
input wire [16-1:0] in);
    wire in0;
    wire in1;
    wire in2;
    wire in3;
    wire in4;
    wire in5;
    wire in6;
    wire in7;
    wire in8;
    wire in9;
    wire in10;
    wire in11;
    wire in12;
    wire in13;
    wire in14;
    wire in15;
    assign in0 = in[0];
    assign in1 = in[1];
    assign in2 = in[2];
    assign in3 = in[3];
    assign in4 = in[4];
    assign in5 = in[5];
    assign in6 = in[6];
    assign in7 = in[7];
    assign in8 = in[8];
    assign in9 = in[9];
    assign in10 = in[10];
    assign in11 = in[11];
    assign in12 = in[12];
    assign in13 = in[13];
    assign in14 = in[14];
    assign in15 = in[15];
    wire in0;
    wire w1;
    wire w20;
    wire w9;
    wire w21;
    wire w17;
    wire w22;
    wire w13;
    wire w23;
    wire w18;
    wire w24;
    wire w16;
    wire w25;
    wire w19;
    wire w26;
    wire w15;
    assign out[0] = in0;
    assign out[1] = w1;
    assign out[2] = w20;
    assign out[3] = w9;
    assign out[4] = w21;
    assign out[5] = w17;
    assign out[6] = w22;
    assign out[7] = w13;
    assign out[8] = w23;
    assign out[9] = w18;
    assign out[10] = w24;
    assign out[11] = w16;
    assign out[12] = w25;
    assign out[13] = w19;
    assign out[14] = w26;
    assign out[15] = w15;
    or or0(w1, in0, in1);
    wire w6;
    or or1(w6, in10, in11);
    wire w7;
    or or2(w7, in12, in13);
    wire w8;
    or or3(w8, in14, in15);
    wire w2;
    or or4(w2, in2, in3);
    wire w3;
    or or5(w3, in4, in5);
    wire w4;
    or or6(w4, in6, in7);
    wire w5;
    or or7(w5, in8, in9);
    or or8(w20, w1, in2);
    or or9(w9, w1, w2);
    wire w10;
    or or10(w10, w3, w4);
    wire w11;
    or or11(w11, w5, w6);
    wire w12;
    or or12(w12, w7, w8);
    wire w14;
    or or13(w14, w11, w12);
    or or14(w21, w9, in4);
    or or15(w13, w9, w10);
    or or16(w17, w9, w3);
    or or17(w23, w13, in8);
    or or18(w16, w13, w11);
    or or19(w15, w13, w14);
    or or20(w18, w13, w5);
    or or21(w22, w17, in6);
    or or22(w25, w16, in12);
    or or23(w19, w16, w7);
    or or24(w24, w18, in10);
    or or25(w26, w19, in14);
endmodule
