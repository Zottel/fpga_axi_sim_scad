`default_nettype none

module top
#(
  parameter integer C_S_AXI_CONTROL_DATA_WIDTH = 32,
  parameter integer C_S_AXI_CONTROL_ADDR_WIDTH = 6,
  parameter integer C_M_AXI_PROGMEM_ID_WIDTH = 1,
  parameter integer C_M_AXI_PROGMEM_DATA_WIDTH = 256,
  parameter integer C_M_AXI_PROGMEM_ADDR_WIDTH = 64,
  parameter integer C_M_AXI_GMEM_ID_WIDTH = 1,
  parameter integer C_M_AXI_GMEM_DATA_WIDTH = 64,
  parameter integer C_M_AXI_GMEM_ADDR_WIDTH = 64
)(
    input wire ap_clk,
    input wire ap_rst_n,
  input wire  s_axi_control_AWVALID,
  input wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_AWADDR,
  input wire  s_axi_control_WVALID,
  input wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_WDATA,
  input wire [C_S_AXI_CONTROL_DATA_WIDTH/8-1:0] s_axi_control_WSTRB,
  input wire  s_axi_control_ARVALID,
  input wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_ARADDR,
  input wire  s_axi_control_RREADY,
  input wire  s_axi_control_BREADY,
  output wire  s_axi_control_AWREADY,
  output wire  s_axi_control_WREADY,
  output wire  s_axi_control_ARREADY,
  output wire  s_axi_control_RVALID,
  output wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_RDATA,
  output wire [1:0] s_axi_control_RRESP,
  output wire  s_axi_control_BVALID,
  output wire [1:0] s_axi_control_BRESP,
  input wire  m_axi_progmem_AWREADY,
  input wire  m_axi_progmem_WREADY,
  input wire  m_axi_progmem_ARREADY,
  input wire  m_axi_progmem_RVALID,
  input wire [C_M_AXI_PROGMEM_DATA_WIDTH-1:0] m_axi_progmem_RDATA,
  input wire  m_axi_progmem_RLAST,
  input wire [C_M_AXI_PROGMEM_ID_WIDTH-1:0] m_axi_progmem_RID,
  input wire [1:0] m_axi_progmem_RRESP,
  input wire  m_axi_progmem_BVALID,
  input wire [C_M_AXI_PROGMEM_ID_WIDTH-1:0] m_axi_progmem_BID,
  input wire [1:0] m_axi_progmem_BRESP,
  output wire  m_axi_progmem_AWVALID,
  output wire [C_M_AXI_PROGMEM_ADDR_WIDTH-1:0] m_axi_progmem_AWADDR,
  output wire [C_M_AXI_PROGMEM_ID_WIDTH-1:0] m_axi_progmem_AWID,
  output wire [7:0] m_axi_progmem_AWLEN,
  output wire [2:0] m_axi_progmem_AWSIZE,
  output wire [1:0] m_axi_progmem_AWBURST,
  output wire [1:0] m_axi_progmem_AWLOCK,
  output wire [3:0] m_axi_progmem_AWCACHE,
  output wire [2:0] m_axi_progmem_AWPROT,
  output wire [3:0] m_axi_progmem_AWQOS,
  output wire [3:0] m_axi_progmem_AWREGION,
  output wire  m_axi_progmem_WVALID,
  output wire [C_M_AXI_PROGMEM_DATA_WIDTH-1:0] m_axi_progmem_WDATA,
  output wire [C_M_AXI_PROGMEM_DATA_WIDTH/8-1:0] m_axi_progmem_WSTRB,
  output wire  m_axi_progmem_WLAST,
  output wire  m_axi_progmem_ARVALID,
  output wire [C_M_AXI_PROGMEM_ADDR_WIDTH-1:0] m_axi_progmem_ARADDR,
  output wire [C_M_AXI_PROGMEM_ID_WIDTH-1:0] m_axi_progmem_ARID,
  output wire [7:0] m_axi_progmem_ARLEN,
  output wire [2:0] m_axi_progmem_ARSIZE,
  output wire [1:0] m_axi_progmem_ARBURST,
  output wire [1:0] m_axi_progmem_ARLOCK,
  output wire [3:0] m_axi_progmem_ARCACHE,
  output wire [2:0] m_axi_progmem_ARPROT,
  output wire [3:0] m_axi_progmem_ARQOS,
  output wire [3:0] m_axi_progmem_ARREGION,
  output wire  m_axi_progmem_RREADY,
  output wire  m_axi_progmem_BREADY,
  input wire  m_axi_gmem_AWREADY,
  input wire  m_axi_gmem_WREADY,
  input wire  m_axi_gmem_ARREADY,
  input wire  m_axi_gmem_RVALID,
  input wire [C_M_AXI_GMEM_DATA_WIDTH-1:0] m_axi_gmem_RDATA,
  input wire  m_axi_gmem_RLAST,
  input wire [C_M_AXI_GMEM_ID_WIDTH-1:0] m_axi_gmem_RID,
  input wire [1:0] m_axi_gmem_RRESP,
  input wire  m_axi_gmem_BVALID,
  input wire [C_M_AXI_GMEM_ID_WIDTH-1:0] m_axi_gmem_BID,
  input wire [1:0] m_axi_gmem_BRESP,
  output wire  m_axi_gmem_AWVALID,
  output wire [C_M_AXI_GMEM_ADDR_WIDTH-1:0] m_axi_gmem_AWADDR,
  output wire [C_M_AXI_GMEM_ID_WIDTH-1:0] m_axi_gmem_AWID,
  output wire [7:0] m_axi_gmem_AWLEN,
  output wire [2:0] m_axi_gmem_AWSIZE,
  output wire [1:0] m_axi_gmem_AWBURST,
  output wire [1:0] m_axi_gmem_AWLOCK,
  output wire [3:0] m_axi_gmem_AWCACHE,
  output wire [2:0] m_axi_gmem_AWPROT,
  output wire [3:0] m_axi_gmem_AWQOS,
  output wire [3:0] m_axi_gmem_AWREGION,
  output wire  m_axi_gmem_WVALID,
  output wire [C_M_AXI_GMEM_DATA_WIDTH-1:0] m_axi_gmem_WDATA,
  output wire [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m_axi_gmem_WSTRB,
  output wire  m_axi_gmem_WLAST,
  output wire  m_axi_gmem_ARVALID,
  output wire [C_M_AXI_GMEM_ADDR_WIDTH-1:0] m_axi_gmem_ARADDR,
  output wire [C_M_AXI_GMEM_ID_WIDTH-1:0] m_axi_gmem_ARID,
  output wire [7:0] m_axi_gmem_ARLEN,
  output wire [2:0] m_axi_gmem_ARSIZE,
  output wire [1:0] m_axi_gmem_ARBURST,
  output wire [1:0] m_axi_gmem_ARLOCK,
  output wire [3:0] m_axi_gmem_ARCACHE,
  output wire [2:0] m_axi_gmem_ARPROT,
  output wire [3:0] m_axi_gmem_ARQOS,
  output wire [3:0] m_axi_gmem_ARREGION,
  output wire  m_axi_gmem_RREADY,
  output wire  m_axi_gmem_BREADY
);
  
  top_int #(
    .C_S_AXI_CONTROL_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH),
    .C_S_AXI_CONTROL_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_M_AXI_PROGMEM_ID_WIDTH(C_M_AXI_PROGMEM_ID_WIDTH),
    .C_M_AXI_PROGMEM_DATA_WIDTH(C_M_AXI_PROGMEM_DATA_WIDTH),
    .C_M_AXI_PROGMEM_ADDR_WIDTH(C_M_AXI_PROGMEM_ADDR_WIDTH),
    .C_M_AXI_GMEM_ID_WIDTH(C_M_AXI_GMEM_ID_WIDTH),
    .C_M_AXI_GMEM_DATA_WIDTH(C_M_AXI_GMEM_DATA_WIDTH),
    .C_M_AXI_GMEM_ADDR_WIDTH(C_M_AXI_GMEM_ADDR_WIDTH)
  ) top_int_inst (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .s_axi_control_AWVALID(s_axi_control_AWVALID),
    .s_axi_control_AWADDR(s_axi_control_AWADDR),
    .s_axi_control_WVALID(s_axi_control_WVALID),
    .s_axi_control_WDATA(s_axi_control_WDATA),
    .s_axi_control_WSTRB(s_axi_control_WSTRB),
    .s_axi_control_ARVALID(s_axi_control_ARVALID),
    .s_axi_control_ARADDR(s_axi_control_ARADDR),
    .s_axi_control_RREADY(s_axi_control_RREADY),
    .s_axi_control_BREADY(s_axi_control_BREADY),
    .s_axi_control_AWREADY(s_axi_control_AWREADY),
    .s_axi_control_WREADY(s_axi_control_WREADY),
    .s_axi_control_ARREADY(s_axi_control_ARREADY),
    .s_axi_control_RVALID(s_axi_control_RVALID),
    .s_axi_control_RDATA(s_axi_control_RDATA),
    .s_axi_control_RRESP(s_axi_control_RRESP),
    .s_axi_control_BVALID(s_axi_control_BVALID),
    .s_axi_control_BRESP(s_axi_control_BRESP),
    .m_axi_progmem_AWREADY(m_axi_progmem_AWREADY),
    .m_axi_progmem_WREADY(m_axi_progmem_WREADY),
    .m_axi_progmem_ARREADY(m_axi_progmem_ARREADY),
    .m_axi_progmem_RVALID(m_axi_progmem_RVALID),
    .m_axi_progmem_RDATA(m_axi_progmem_RDATA),
    .m_axi_progmem_RLAST(m_axi_progmem_RLAST),
    .m_axi_progmem_RID(m_axi_progmem_RID),
    .m_axi_progmem_RRESP(m_axi_progmem_RRESP),
    .m_axi_progmem_BVALID(m_axi_progmem_BVALID),
    .m_axi_progmem_BID(m_axi_progmem_BID),
    .m_axi_progmem_BRESP(m_axi_progmem_BRESP),
    .m_axi_progmem_AWVALID(m_axi_progmem_AWVALID),
    .m_axi_progmem_AWADDR(m_axi_progmem_AWADDR),
    .m_axi_progmem_AWID(m_axi_progmem_AWID),
    .m_axi_progmem_AWLEN(m_axi_progmem_AWLEN),
    .m_axi_progmem_AWSIZE(m_axi_progmem_AWSIZE),
    .m_axi_progmem_AWBURST(m_axi_progmem_AWBURST),
    .m_axi_progmem_AWLOCK(m_axi_progmem_AWLOCK),
    .m_axi_progmem_AWCACHE(m_axi_progmem_AWCACHE),
    .m_axi_progmem_AWPROT(m_axi_progmem_AWPROT),
    .m_axi_progmem_AWQOS(m_axi_progmem_AWQOS),
    .m_axi_progmem_AWREGION(m_axi_progmem_AWREGION),
    .m_axi_progmem_WVALID(m_axi_progmem_WVALID),
    .m_axi_progmem_WDATA(m_axi_progmem_WDATA),
    .m_axi_progmem_WSTRB(m_axi_progmem_WSTRB),
    .m_axi_progmem_WLAST(m_axi_progmem_WLAST),
    .m_axi_progmem_ARVALID(m_axi_progmem_ARVALID),
    .m_axi_progmem_ARADDR(m_axi_progmem_ARADDR),
    .m_axi_progmem_ARID(m_axi_progmem_ARID),
    .m_axi_progmem_ARLEN(m_axi_progmem_ARLEN),
    .m_axi_progmem_ARSIZE(m_axi_progmem_ARSIZE),
    .m_axi_progmem_ARBURST(m_axi_progmem_ARBURST),
    .m_axi_progmem_ARLOCK(m_axi_progmem_ARLOCK),
    .m_axi_progmem_ARCACHE(m_axi_progmem_ARCACHE),
    .m_axi_progmem_ARPROT(m_axi_progmem_ARPROT),
    .m_axi_progmem_ARQOS(m_axi_progmem_ARQOS),
    .m_axi_progmem_ARREGION(m_axi_progmem_ARREGION),
    .m_axi_progmem_RREADY(m_axi_progmem_RREADY),
    .m_axi_progmem_BREADY(m_axi_progmem_BREADY),
    .m_axi_gmem_AWREADY(m_axi_gmem_AWREADY),
    .m_axi_gmem_WREADY(m_axi_gmem_WREADY),
    .m_axi_gmem_ARREADY(m_axi_gmem_ARREADY),
    .m_axi_gmem_RVALID(m_axi_gmem_RVALID),
    .m_axi_gmem_RDATA(m_axi_gmem_RDATA),
    .m_axi_gmem_RLAST(m_axi_gmem_RLAST),
    .m_axi_gmem_RID(m_axi_gmem_RID),
    .m_axi_gmem_RRESP(m_axi_gmem_RRESP),
    .m_axi_gmem_BVALID(m_axi_gmem_BVALID),
    .m_axi_gmem_BID(m_axi_gmem_BID),
    .m_axi_gmem_BRESP(m_axi_gmem_BRESP),
    .m_axi_gmem_AWVALID(m_axi_gmem_AWVALID),
    .m_axi_gmem_AWADDR(m_axi_gmem_AWADDR),
    .m_axi_gmem_AWID(m_axi_gmem_AWID),
    .m_axi_gmem_AWLEN(m_axi_gmem_AWLEN),
    .m_axi_gmem_AWSIZE(m_axi_gmem_AWSIZE),
    .m_axi_gmem_AWBURST(m_axi_gmem_AWBURST),
    .m_axi_gmem_AWLOCK(m_axi_gmem_AWLOCK),
    .m_axi_gmem_AWCACHE(m_axi_gmem_AWCACHE),
    .m_axi_gmem_AWPROT(m_axi_gmem_AWPROT),
    .m_axi_gmem_AWQOS(m_axi_gmem_AWQOS),
    .m_axi_gmem_AWREGION(m_axi_gmem_AWREGION),
    .m_axi_gmem_WVALID(m_axi_gmem_WVALID),
    .m_axi_gmem_WDATA(m_axi_gmem_WDATA),
    .m_axi_gmem_WSTRB(m_axi_gmem_WSTRB),
    .m_axi_gmem_WLAST(m_axi_gmem_WLAST),
    .m_axi_gmem_ARVALID(m_axi_gmem_ARVALID),
    .m_axi_gmem_ARADDR(m_axi_gmem_ARADDR),
    .m_axi_gmem_ARID(m_axi_gmem_ARID),
    .m_axi_gmem_ARLEN(m_axi_gmem_ARLEN),
    .m_axi_gmem_ARSIZE(m_axi_gmem_ARSIZE),
    .m_axi_gmem_ARBURST(m_axi_gmem_ARBURST),
    .m_axi_gmem_ARLOCK(m_axi_gmem_ARLOCK),
    .m_axi_gmem_ARCACHE(m_axi_gmem_ARCACHE),
    .m_axi_gmem_ARPROT(m_axi_gmem_ARPROT),
    .m_axi_gmem_ARQOS(m_axi_gmem_ARQOS),
    .m_axi_gmem_ARREGION(m_axi_gmem_ARREGION),
    .m_axi_gmem_RREADY(m_axi_gmem_RREADY),
    .m_axi_gmem_BREADY(m_axi_gmem_BREADY)
  );  
endmodule
